-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2016.12.27910

-- Build Date:         Dec 21 2016 18:07:02

-- File Generated:     Apr 1 2017 16:19:35

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "uart_rx_fsm" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of uart_rx_fsm
entity uart_rx_fsm is
port (
    i_no_of_data_bits : in std_logic_vector(1 downto 0);
    o_rx_data : out std_logic_vector(7 downto 0);
    i_start_rx : in std_logic;
    o_parity_error : out std_logic;
    i_clear_linestatusreg : in std_logic;
    o_rx_data_ready : out std_logic;
    i_stick_parity_en : in std_logic;
    i_rx_clk : in std_logic;
    i_clear_rxdataready : in std_logic;
    o_timeout : out std_logic;
    o_framing_error : out std_logic;
    i_serial_data : in std_logic;
    i_parity_even : in std_logic;
    i_parity_en : in std_logic;
    i_int_serial_data : in std_logic;
    i_clk : in std_logic;
    o_break_interrupt : out std_logic;
    i_rst : in std_logic;
    bit_sample_en : out std_logic;
    i_loopback_en : in std_logic);
end uart_rx_fsm;

-- Architecture of uart_rx_fsm
-- View name is \INTERFACE\
architecture \INTERFACE\ of uart_rx_fsm is

signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1992\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1959\ : std_logic;
signal \N__1956\ : std_logic;
signal \N__1953\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal i_rst_ibuf_gb_io_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal o_rx_data_c_6 : std_logic;
signal o_rx_data_c_7 : std_logic;
signal o_rx_data_c_1 : std_logic;
signal o_rx_data_c_2 : std_logic;
signal o_rx_data_c_0 : std_logic;
signal o_rx_data_c_4 : std_logic;
signal i_serial_data_c : std_logic;
signal i_loopback_en_c : std_logic;
signal i_int_serial_data_c : std_logic;
signal state_ns_i_i_a2_0_9 : std_logic;
signal o_rx_data_c_3 : std_logic;
signal o_rx_data_c_5 : std_logic;
signal \N_187\ : std_logic;
signal \N_176_cascade_\ : std_logic;
signal \N_176\ : std_logic;
signal rx_data_35_0_iv_0_a2_0_1_3 : std_logic;
signal \N_148_cascade_\ : std_logic;
signal rx_data_35_0_iv_0_a2_0_1_5 : std_logic;
signal \N_152_cascade_\ : std_logic;
signal \N_157_cascade_\ : std_logic;
signal rx_data_35_0_iv_0_a2_3_out_0 : std_logic;
signal rx_data_35_0_iv_0_a2_0_1_s_0_7 : std_logic;
signal \rx_data_35_0_iv_0_a2_0_1_s_0_7_cascade_\ : std_logic;
signal \N_183_cascade_\ : std_logic;
signal rx_data_35_0_iv_0_a2_0_1_s_0_0_9 : std_logic;
signal \rx_data_35_0_iv_0_a2_0_1_s_0_0_9_cascade_\ : std_logic;
signal \state_ns_i_i_0_a2_0_8_cascade_\ : std_logic;
signal \rx_data_35_0_iv_0_a2_0_0_4_cascade_\ : std_logic;
signal i_no_of_data_bits_c_1 : std_logic;
signal \stateZ0Z_8\ : std_logic;
signal \state_fastZ0Z_6\ : std_logic;
signal \stateZ0Z_6\ : std_logic;
signal \N_378\ : std_logic;
signal \data_validationZ0\ : std_logic;
signal break_interrupt_e_sn : std_logic;
signal break_interrupt_e_rn_0 : std_logic;
signal \break_interrupt_0_sqmuxa_0_a2_6_cascade_\ : std_logic;
signal break_interrupt_0_sqmuxa_0_a2_7 : std_logic;
signal \un1_rx_data_0_sqmuxa_2_i_a2_d_0_0_cascade_\ : std_logic;
signal un1_framing_error_0_sqmuxa_0_i : std_logic;
signal \N_13_i_1_1_cascade_\ : std_logic;
signal \clear_data_readyZ0\ : std_logic;
signal \N_386\ : std_logic;
signal \N_13_i_1\ : std_logic;
signal \N_165_cascade_\ : std_logic;
signal rx_data_35_0_iv_0_a2_1_0_0 : std_logic;
signal \N_143_cascade_\ : std_logic;
signal \rx_dataZ0Z_0\ : std_logic;
signal \N_115\ : std_logic;
signal \N_174\ : std_logic;
signal \N_150_cascade_\ : std_logic;
signal rx_data_35_0_iv_0_a2_0_1_4 : std_logic;
signal \N_142_cascade_\ : std_logic;
signal \N_155\ : std_logic;
signal \rx_data_RNO_2Z0Z_1_cascade_\ : std_logic;
signal \rx_data_RNO_1Z0Z_1_cascade_\ : std_logic;
signal rx_data_35_0_i_1_1 : std_logic;
signal \N_92_cascade_\ : std_logic;
signal \N_183\ : std_logic;
signal \N_147_cascade_\ : std_logic;
signal \stateZ0Z_9\ : std_logic;
signal \N_182\ : std_logic;
signal \modem_serial_data_repZ0Z1\ : std_logic;
signal \N_377\ : std_logic;
signal \rx_sampling_clock_reg2_fastZ0\ : std_logic;
signal \stateZ0Z_5\ : std_logic;
signal \stateZ0Z_4\ : std_logic;
signal \stateZ0Z_3\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal timeout_counter_cry_0 : std_logic;
signal timeout_counter_cry_1 : std_logic;
signal timeout_counter_cry_2 : std_logic;
signal timeout_counter_cry_3 : std_logic;
signal timeout_counter_cry_4 : std_logic;
signal \o_timeout5_3_cascade_\ : std_logic;
signal o_timeout_c : std_logic;
signal \timeout_counterZ0Z_0\ : std_logic;
signal \timeout_counterZ0Z_1\ : std_logic;
signal \timeout_counterZ0Z_2\ : std_logic;
signal \timeout_counterZ0Z_3\ : std_logic;
signal \o2_cascade_\ : std_logic;
signal \timeout_counter_RNI09R61Z0Z_5\ : std_logic;
signal i_clear_rxdataready_c : std_logic;
signal timeout_counter_s_4 : std_logic;
signal \timeout_counterZ0Z_4\ : std_logic;
signal \clearrxdatareadyZ0Z1\ : std_logic;
signal \N_345_0_i\ : std_logic;
signal timeout_counter_s_5 : std_logic;
signal \timeout_counterZ0Z_5\ : std_logic;
signal timeout_countere_0_i : std_logic;
signal o_break_interrupt_c : std_logic;
signal o_parity_error_c : std_logic;
signal \rx_data_ready_regZ0Z1\ : std_logic;
signal \rx_data_ready_regZ0Z2\ : std_logic;
signal o_rx_data_ready_c : std_logic;
signal i_no_of_data_bits_c_0 : std_logic;
signal \stateZ0Z_7\ : std_logic;
signal \N_181\ : std_logic;
signal \rx_sampling_clock_regZ0Z1\ : std_logic;
signal \stateZ0Z_2\ : std_logic;
signal \N_380_cascade_\ : std_logic;
signal \N_161\ : std_logic;
signal \N_379\ : std_logic;
signal \N_142\ : std_logic;
signal \N_159\ : std_logic;
signal \N_16_i\ : std_logic;
signal \rx_sampling_clock_regZ0Z2\ : std_logic;
signal \modem_serial_data_fastZ0\ : std_logic;
signal \N_88\ : std_logic;
signal \rx_sampling_startZ0\ : std_logic;
signal \N_103_cascade_\ : std_logic;
signal timeout_counter_2_sqmuxa : std_logic;
signal \rx_sampling_counterZ0Z_2\ : std_logic;
signal \rx_sampling_counterZ0Z_1\ : std_logic;
signal \rx_sampling_counter_RNO_0Z0Z_3\ : std_logic;
signal \rx_sampling_counterZ0Z_0\ : std_logic;
signal \rx_sampling_counterZ0Z_3\ : std_logic;
signal i_rx_clk_c_g : std_logic;
signal i_clear_linestatusreg_c : std_logic;
signal i_start_rx_c : std_logic;
signal \stateZ0Z_0\ : std_logic;
signal \timeout_counter_beginZ0\ : std_logic;
signal \N_42\ : std_logic;
signal i_rx_clk_c : std_logic;
signal \rx_sampling_clockZ0\ : std_logic;
signal \rx_sampling_clock_reg1_fastZ0\ : std_logic;
signal \stateZ0Z_10\ : std_logic;
signal \rx_clk_regZ0Z1\ : std_logic;
signal \rx_clk_regZ0Z2\ : std_logic;
signal o_framing_error_c : std_logic;
signal \clear_line_statusZ0\ : std_logic;
signal i_parity_en_c : std_logic;
signal i_stick_parity_en_c : std_logic;
signal \stick_parity_bitZ0\ : std_logic;
signal \rx_dataZ0Z_3\ : std_logic;
signal \rx_dataZ0Z_4\ : std_logic;
signal \rx_dataZ0Z_5\ : std_logic;
signal \rx_dataZ0Z_2\ : std_logic;
signal \N_103\ : std_logic;
signal \N_103_0\ : std_logic;
signal \rx_dataZ0Z_8\ : std_logic;
signal \rx_dataZ0Z_7\ : std_logic;
signal \rx_dataZ0Z_9\ : std_logic;
signal \rx_dataZ0Z_1\ : std_logic;
signal parity_error_e_1 : std_logic;
signal i_parity_even_c : std_logic;
signal \N_398\ : std_logic;
signal \parity_errorZ0\ : std_logic;
signal \N_18_i_1\ : std_logic;
signal check_bit_3_1 : std_logic;
signal check_bit_2_5 : std_logic;
signal \rx_dataZ0Z_6\ : std_logic;
signal \stateZ0Z_11\ : std_logic;
signal \check_bitZ0\ : std_logic;
signal \modem_serial_dataZ0\ : std_logic;
signal \stateZ0Z_1\ : std_logic;
signal \framing_errorZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal i_clk_c_g : std_logic;
signal un1_rx_data_0_sqmuxa_1_0_i : std_logic;
signal i_rst_c_g : std_logic;

signal i_clk_wire : std_logic;
signal o_rx_data_wire : std_logic_vector(7 downto 0);
signal o_framing_error_wire : std_logic;
signal i_start_rx_wire : std_logic;
signal o_break_interrupt_wire : std_logic;
signal i_int_serial_data_wire : std_logic;
signal i_parity_en_wire : std_logic;
signal bit_sample_en_wire : std_logic;
signal i_no_of_data_bits_wire : std_logic_vector(1 downto 0);
signal i_rx_clk_wire : std_logic;
signal i_clear_rxdataready_wire : std_logic;
signal o_timeout_wire : std_logic;
signal i_stick_parity_en_wire : std_logic;
signal i_loopback_en_wire : std_logic;
signal i_clear_linestatusreg_wire : std_logic;
signal o_rx_data_ready_wire : std_logic;
signal o_parity_error_wire : std_logic;
signal i_serial_data_wire : std_logic;
signal i_parity_even_wire : std_logic;
signal i_rst_wire : std_logic;

begin
    i_clk_wire <= i_clk;
    o_rx_data <= o_rx_data_wire;
    o_framing_error <= o_framing_error_wire;
    i_start_rx_wire <= i_start_rx;
    o_break_interrupt <= o_break_interrupt_wire;
    i_int_serial_data_wire <= i_int_serial_data;
    i_parity_en_wire <= i_parity_en;
    bit_sample_en <= bit_sample_en_wire;
    i_no_of_data_bits_wire <= i_no_of_data_bits;
    i_rx_clk_wire <= i_rx_clk;
    i_clear_rxdataready_wire <= i_clear_rxdataready;
    o_timeout <= o_timeout_wire;
    i_stick_parity_en_wire <= i_stick_parity_en;
    i_loopback_en_wire <= i_loopback_en;
    i_clear_linestatusreg_wire <= i_clear_linestatusreg;
    o_rx_data_ready <= o_rx_data_ready_wire;
    o_parity_error <= o_parity_error_wire;
    i_serial_data_wire <= i_serial_data;
    i_parity_even_wire <= i_parity_even;
    i_rst_wire <= i_rst;

    \i_clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5578\,
            GLOBALBUFFEROUTPUT => i_clk_c_g
        );

    \i_clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5580\,
            DIN => \N__5579\,
            DOUT => \N__5578\,
            PACKAGEPIN => i_clk_wire
        );

    \i_clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5580\,
            PADOUT => \N__5579\,
            PADIN => \N__5578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5569\,
            DIN => \N__5568\,
            DOUT => \N__5567\,
            PACKAGEPIN => o_rx_data_wire(5)
        );

    \o_rx_data_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5569\,
            PADOUT => \N__5568\,
            PADIN => \N__5567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_framing_error_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5560\,
            DIN => \N__5559\,
            DOUT => \N__5558\,
            PACKAGEPIN => o_framing_error_wire
        );

    \o_framing_error_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5560\,
            PADOUT => \N__5559\,
            PADIN => \N__5558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4344\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_start_rx_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5551\,
            DIN => \N__5550\,
            DOUT => \N__5549\,
            PACKAGEPIN => i_start_rx_wire
        );

    \i_start_rx_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5551\,
            PADOUT => \N__5550\,
            PADIN => \N__5549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_start_rx_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_break_interrupt_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5542\,
            DIN => \N__5541\,
            DOUT => \N__5540\,
            PACKAGEPIN => o_break_interrupt_wire
        );

    \o_break_interrupt_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5542\,
            PADOUT => \N__5541\,
            PADIN => \N__5540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3858\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5533\,
            DIN => \N__5532\,
            DOUT => \N__5531\,
            PACKAGEPIN => o_rx_data_wire(2)
        );

    \o_rx_data_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5533\,
            PADOUT => \N__5532\,
            PADIN => \N__5531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1998\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5524\,
            DIN => \N__5523\,
            DOUT => \N__5522\,
            PACKAGEPIN => o_rx_data_wire(7)
        );

    \o_rx_data_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5524\,
            PADOUT => \N__5523\,
            PADIN => \N__5522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_int_serial_data_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5515\,
            DIN => \N__5514\,
            DOUT => \N__5513\,
            PACKAGEPIN => i_int_serial_data_wire
        );

    \i_int_serial_data_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5515\,
            PADOUT => \N__5514\,
            PADIN => \N__5513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_int_serial_data_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_parity_en_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5506\,
            DIN => \N__5505\,
            DOUT => \N__5504\,
            PACKAGEPIN => i_parity_en_wire
        );

    \i_parity_en_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5506\,
            PADOUT => \N__5505\,
            PADIN => \N__5504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_parity_en_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \bit_sample_en_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5497\,
            DIN => \N__5496\,
            DOUT => \N__5495\,
            PACKAGEPIN => bit_sample_en_wire
        );

    \bit_sample_en_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5497\,
            PADOUT => \N__5496\,
            PADIN => \N__5495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5133\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_no_of_data_bits_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5488\,
            DIN => \N__5487\,
            DOUT => \N__5486\,
            PACKAGEPIN => i_no_of_data_bits_wire(0)
        );

    \i_no_of_data_bits_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5488\,
            PADOUT => \N__5487\,
            PADIN => \N__5486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_no_of_data_bits_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_rx_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5479\,
            DIN => \N__5478\,
            DOUT => \N__5477\,
            PACKAGEPIN => i_rx_clk_wire
        );

    \i_rx_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5479\,
            PADOUT => \N__5478\,
            PADIN => \N__5477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_rx_clk_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_clear_rxdataready_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5470\,
            DIN => \N__5469\,
            DOUT => \N__5468\,
            PACKAGEPIN => i_clear_rxdataready_wire
        );

    \i_clear_rxdataready_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5470\,
            PADOUT => \N__5469\,
            PADIN => \N__5468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_clear_rxdataready_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_timeout_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5461\,
            DIN => \N__5460\,
            DOUT => \N__5459\,
            PACKAGEPIN => o_timeout_wire
        );

    \o_timeout_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5461\,
            PADOUT => \N__5460\,
            PADIN => \N__5459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5452\,
            DIN => \N__5451\,
            DOUT => \N__5450\,
            PACKAGEPIN => o_rx_data_wire(4)
        );

    \o_rx_data_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5452\,
            PADOUT => \N__5451\,
            PADIN => \N__5450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1971\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_no_of_data_bits_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5443\,
            DIN => \N__5442\,
            DOUT => \N__5441\,
            PACKAGEPIN => i_no_of_data_bits_wire(1)
        );

    \i_no_of_data_bits_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5443\,
            PADOUT => \N__5442\,
            PADIN => \N__5441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_no_of_data_bits_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_stick_parity_en_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5434\,
            DIN => \N__5433\,
            DOUT => \N__5432\,
            PACKAGEPIN => i_stick_parity_en_wire
        );

    \i_stick_parity_en_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5434\,
            PADOUT => \N__5433\,
            PADIN => \N__5432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_stick_parity_en_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5425\,
            DIN => \N__5424\,
            DOUT => \N__5423\,
            PACKAGEPIN => o_rx_data_wire(0)
        );

    \o_rx_data_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5425\,
            PADOUT => \N__5424\,
            PADIN => \N__5423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1986\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_loopback_en_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5416\,
            DIN => \N__5415\,
            DOUT => \N__5414\,
            PACKAGEPIN => i_loopback_en_wire
        );

    \i_loopback_en_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5416\,
            PADOUT => \N__5415\,
            PADIN => \N__5414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_loopback_en_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5407\,
            DIN => \N__5406\,
            DOUT => \N__5405\,
            PACKAGEPIN => o_rx_data_wire(1)
        );

    \o_rx_data_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5407\,
            PADOUT => \N__5406\,
            PADIN => \N__5405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2013\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_clear_linestatusreg_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5398\,
            DIN => \N__5397\,
            DOUT => \N__5396\,
            PACKAGEPIN => i_clear_linestatusreg_wire
        );

    \i_clear_linestatusreg_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5398\,
            PADOUT => \N__5397\,
            PADIN => \N__5396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_clear_linestatusreg_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5389\,
            DIN => \N__5388\,
            DOUT => \N__5387\,
            PACKAGEPIN => o_rx_data_wire(6)
        );

    \o_rx_data_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5389\,
            PADOUT => \N__5388\,
            PADIN => \N__5387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_ready_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5380\,
            DIN => \N__5379\,
            DOUT => \N__5378\,
            PACKAGEPIN => o_rx_data_ready_wire
        );

    \o_rx_data_ready_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5380\,
            PADOUT => \N__5379\,
            PADIN => \N__5378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3786\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_parity_error_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5371\,
            DIN => \N__5370\,
            DOUT => \N__5369\,
            PACKAGEPIN => o_parity_error_wire
        );

    \o_parity_error_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5371\,
            PADOUT => \N__5370\,
            PADIN => \N__5369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_rx_data_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5362\,
            DIN => \N__5361\,
            DOUT => \N__5360\,
            PACKAGEPIN => o_rx_data_wire(3)
        );

    \o_rx_data_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5362\,
            PADOUT => \N__5361\,
            PADIN => \N__5360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2061\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_serial_data_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5353\,
            DIN => \N__5352\,
            DOUT => \N__5351\,
            PACKAGEPIN => i_serial_data_wire
        );

    \i_serial_data_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5353\,
            PADOUT => \N__5352\,
            PADIN => \N__5351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_serial_data_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_parity_even_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5344\,
            DIN => \N__5343\,
            DOUT => \N__5342\,
            PACKAGEPIN => i_parity_even_wire
        );

    \i_parity_even_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5344\,
            PADOUT => \N__5343\,
            PADIN => \N__5342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_parity_even_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_rst_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5335\,
            DIN => \N__5334\,
            DOUT => \N__5333\,
            PACKAGEPIN => i_rst_wire
        );

    \i_rst_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5335\,
            PADOUT => \N__5334\,
            PADIN => \N__5333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_rst_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1290\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5312\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5309\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5312\,
            I => \N__5305\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5309\,
            I => \N__5302\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5298\
        );

    \I__1285\ : Span4Mux_s3_h
    port map (
            O => \N__5305\,
            I => \N__5295\
        );

    \I__1284\ : Span4Mux_s3_h
    port map (
            O => \N__5302\,
            I => \N__5292\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5289\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5298\,
            I => \rx_dataZ0Z_8\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__5295\,
            I => \rx_dataZ0Z_8\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__5292\,
            I => \rx_dataZ0Z_8\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5289\,
            I => \rx_dataZ0Z_8\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5275\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5272\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5269\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5275\,
            I => \N__5263\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5272\,
            I => \N__5263\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5260\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5257\
        );

    \I__1271\ : Span4Mux_v
    port map (
            O => \N__5263\,
            I => \N__5254\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5260\,
            I => \N__5251\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5257\,
            I => \rx_dataZ0Z_7\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__5254\,
            I => \rx_dataZ0Z_7\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__5251\,
            I => \rx_dataZ0Z_7\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5240\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__5243\,
            I => \N__5237\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5234\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5231\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__5234\,
            I => \N__5224\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5224\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__5230\,
            I => \N__5221\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5218\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__5224\,
            I => \N__5215\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5212\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5218\,
            I => \rx_dataZ0Z_9\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__5215\,
            I => \rx_dataZ0Z_9\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5212\,
            I => \rx_dataZ0Z_9\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5201\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__5204\,
            I => \N__5196\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5193\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5190\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5185\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5185\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__5193\,
            I => \N__5182\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5179\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5185\,
            I => \rx_dataZ0Z_1\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__5182\,
            I => \rx_dataZ0Z_1\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__5179\,
            I => \rx_dataZ0Z_1\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5169\,
            I => parity_error_e_1
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__1237\ : Odrv12
    port map (
            O => \N__5157\,
            I => i_parity_even_c
        );

    \I__1236\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5151\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N_398\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5145\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5145\,
            I => \N__5141\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5138\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__5141\,
            I => \parity_errorZ0\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5138\,
            I => \parity_errorZ0\
        );

    \I__1229\ : IoInMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5126\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5121\
        );

    \I__1226\ : IoSpan4Mux
    port map (
            O => \N__5126\,
            I => \N__5118\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__5125\,
            I => \N__5114\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5107\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5121\,
            I => \N__5100\
        );

    \I__1222\ : Span4Mux_s1_h
    port map (
            O => \N__5118\,
            I => \N__5094\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5091\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5088\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__5113\,
            I => \N__5083\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5080\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5077\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__5110\,
            I => \N__5073\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5107\,
            I => \N__5069\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5066\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5063\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5058\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5058\
        );

    \I__1210\ : Span4Mux_s1_h
    port map (
            O => \N__5100\,
            I => \N__5055\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5050\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5050\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5047\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__5094\,
            I => \N__5040\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5040\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5040\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5033\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5033\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5033\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5080\,
            I => \N__5028\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5077\,
            I => \N__5028\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5021\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5021\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5021\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__5069\,
            I => \N_18_i_1\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5066\,
            I => \N_18_i_1\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5063\,
            I => \N_18_i_1\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N_18_i_1\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__5055\,
            I => \N_18_i_1\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5050\,
            I => \N_18_i_1\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N_18_i_1\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__5040\,
            I => \N_18_i_1\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5033\,
            I => \N_18_i_1\
        );

    \I__1186\ : Odrv12
    port map (
            O => \N__5028\,
            I => \N_18_i_1\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N_18_i_1\
        );

    \I__1184\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__4995\,
            I => check_bit_3_1
        );

    \I__1182\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4989\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__4989\,
            I => check_bit_2_5
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__4986\,
            I => \N__4981\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__4985\,
            I => \N__4978\
        );

    \I__1178\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4975\
        );

    \I__1177\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4972\
        );

    \I__1176\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4968\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__4975\,
            I => \N__4963\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4963\
        );

    \I__1173\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4960\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4957\
        );

    \I__1171\ : Span4Mux_s2_h
    port map (
            O => \N__4963\,
            I => \N__4954\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__4960\,
            I => \rx_dataZ0Z_6\
        );

    \I__1169\ : Odrv12
    port map (
            O => \N__4957\,
            I => \rx_dataZ0Z_6\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__4954\,
            I => \rx_dataZ0Z_6\
        );

    \I__1167\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4943\
        );

    \I__1166\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4940\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__4943\,
            I => \N__4934\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4931\
        );

    \I__1163\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4928\
        );

    \I__1162\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4921\
        );

    \I__1161\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4918\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__4934\,
            I => \N__4911\
        );

    \I__1159\ : Span4Mux_v
    port map (
            O => \N__4931\,
            I => \N__4911\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4911\
        );

    \I__1157\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4905\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__4926\,
            I => \N__4901\
        );

    \I__1155\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4898\
        );

    \I__1154\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4895\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__4921\,
            I => \N__4890\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__4918\,
            I => \N__4890\
        );

    \I__1151\ : Span4Mux_h
    port map (
            O => \N__4911\,
            I => \N__4887\
        );

    \I__1150\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4882\
        );

    \I__1149\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4882\
        );

    \I__1148\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4879\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__4905\,
            I => \N__4876\
        );

    \I__1146\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4873\
        );

    \I__1145\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4870\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__4898\,
            I => \stateZ0Z_11\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__4895\,
            I => \stateZ0Z_11\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__4890\,
            I => \stateZ0Z_11\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__4887\,
            I => \stateZ0Z_11\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__4882\,
            I => \stateZ0Z_11\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__4879\,
            I => \stateZ0Z_11\
        );

    \I__1138\ : Odrv12
    port map (
            O => \N__4876\,
            I => \stateZ0Z_11\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__4873\,
            I => \stateZ0Z_11\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__4870\,
            I => \stateZ0Z_11\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__4848\,
            I => \check_bitZ0\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \N__4840\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \N__4837\
        );

    \I__1131\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4833\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4830\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4827\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__4836\,
            I => \N__4822\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__4833\,
            I => \N__4819\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4814\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4827\,
            I => \N__4814\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__4826\,
            I => \N__4811\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__4825\,
            I => \N__4808\
        );

    \I__1122\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4805\
        );

    \I__1121\ : Span4Mux_h
    port map (
            O => \N__4819\,
            I => \N__4800\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__4814\,
            I => \N__4800\
        );

    \I__1119\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4797\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4794\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4787\
        );

    \I__1116\ : Span4Mux_h
    port map (
            O => \N__4800\,
            I => \N__4782\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4782\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4779\
        );

    \I__1113\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4770\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4770\
        );

    \I__1111\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4770\
        );

    \I__1110\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4770\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__4787\,
            I => \N__4767\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__4782\,
            I => \N__4764\
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__4779\,
            I => \modem_serial_dataZ0\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__4770\,
            I => \modem_serial_dataZ0\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__4767\,
            I => \modem_serial_dataZ0\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__4764\,
            I => \modem_serial_dataZ0\
        );

    \I__1103\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4751\
        );

    \I__1102\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4747\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__4751\,
            I => \N__4742\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4739\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4736\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__4746\,
            I => \N__4732\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__4745\,
            I => \N__4729\
        );

    \I__1096\ : Span4Mux_s1_h
    port map (
            O => \N__4742\,
            I => \N__4723\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__4739\,
            I => \N__4720\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__4736\,
            I => \N__4717\
        );

    \I__1093\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4714\
        );

    \I__1092\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4703\
        );

    \I__1091\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4703\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4703\
        );

    \I__1089\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4703\
        );

    \I__1088\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4703\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__4723\,
            I => \stateZ0Z_1\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__4720\,
            I => \stateZ0Z_1\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__4717\,
            I => \stateZ0Z_1\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__4714\,
            I => \stateZ0Z_1\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__4703\,
            I => \stateZ0Z_1\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__4686\,
            I => \N__4683\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__4683\,
            I => \framing_errorZ0\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__4680\,
            I => \N__4608\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__4679\,
            I => \N__4608\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__4678\,
            I => \N__4608\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__4677\,
            I => \N__4608\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__4676\,
            I => \N__4608\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__4675\,
            I => \N__4608\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__4674\,
            I => \N__4608\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__4673\,
            I => \N__4608\
        );

    \I__1070\ : ClkMux
    port map (
            O => \N__4672\,
            I => \N__4608\
        );

    \I__1069\ : ClkMux
    port map (
            O => \N__4671\,
            I => \N__4608\
        );

    \I__1068\ : ClkMux
    port map (
            O => \N__4670\,
            I => \N__4608\
        );

    \I__1067\ : ClkMux
    port map (
            O => \N__4669\,
            I => \N__4608\
        );

    \I__1066\ : ClkMux
    port map (
            O => \N__4668\,
            I => \N__4608\
        );

    \I__1065\ : ClkMux
    port map (
            O => \N__4667\,
            I => \N__4608\
        );

    \I__1064\ : ClkMux
    port map (
            O => \N__4666\,
            I => \N__4608\
        );

    \I__1063\ : ClkMux
    port map (
            O => \N__4665\,
            I => \N__4608\
        );

    \I__1062\ : ClkMux
    port map (
            O => \N__4664\,
            I => \N__4608\
        );

    \I__1061\ : ClkMux
    port map (
            O => \N__4663\,
            I => \N__4608\
        );

    \I__1060\ : ClkMux
    port map (
            O => \N__4662\,
            I => \N__4608\
        );

    \I__1059\ : ClkMux
    port map (
            O => \N__4661\,
            I => \N__4608\
        );

    \I__1058\ : ClkMux
    port map (
            O => \N__4660\,
            I => \N__4608\
        );

    \I__1057\ : ClkMux
    port map (
            O => \N__4659\,
            I => \N__4608\
        );

    \I__1056\ : ClkMux
    port map (
            O => \N__4658\,
            I => \N__4608\
        );

    \I__1055\ : ClkMux
    port map (
            O => \N__4657\,
            I => \N__4608\
        );

    \I__1054\ : GlobalMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__1053\ : gio2CtrlBuf
    port map (
            O => \N__4605\,
            I => i_clk_c_g
        );

    \I__1052\ : CEMux
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__4593\,
            I => un1_rx_data_0_sqmuxa_1_0_i
        );

    \I__1048\ : SRMux
    port map (
            O => \N__4590\,
            I => \N__4512\
        );

    \I__1047\ : SRMux
    port map (
            O => \N__4589\,
            I => \N__4512\
        );

    \I__1046\ : SRMux
    port map (
            O => \N__4588\,
            I => \N__4512\
        );

    \I__1045\ : SRMux
    port map (
            O => \N__4587\,
            I => \N__4512\
        );

    \I__1044\ : SRMux
    port map (
            O => \N__4586\,
            I => \N__4512\
        );

    \I__1043\ : SRMux
    port map (
            O => \N__4585\,
            I => \N__4512\
        );

    \I__1042\ : SRMux
    port map (
            O => \N__4584\,
            I => \N__4512\
        );

    \I__1041\ : SRMux
    port map (
            O => \N__4583\,
            I => \N__4512\
        );

    \I__1040\ : SRMux
    port map (
            O => \N__4582\,
            I => \N__4512\
        );

    \I__1039\ : SRMux
    port map (
            O => \N__4581\,
            I => \N__4512\
        );

    \I__1038\ : SRMux
    port map (
            O => \N__4580\,
            I => \N__4512\
        );

    \I__1037\ : SRMux
    port map (
            O => \N__4579\,
            I => \N__4512\
        );

    \I__1036\ : SRMux
    port map (
            O => \N__4578\,
            I => \N__4512\
        );

    \I__1035\ : SRMux
    port map (
            O => \N__4577\,
            I => \N__4512\
        );

    \I__1034\ : SRMux
    port map (
            O => \N__4576\,
            I => \N__4512\
        );

    \I__1033\ : SRMux
    port map (
            O => \N__4575\,
            I => \N__4512\
        );

    \I__1032\ : SRMux
    port map (
            O => \N__4574\,
            I => \N__4512\
        );

    \I__1031\ : SRMux
    port map (
            O => \N__4573\,
            I => \N__4512\
        );

    \I__1030\ : SRMux
    port map (
            O => \N__4572\,
            I => \N__4512\
        );

    \I__1029\ : SRMux
    port map (
            O => \N__4571\,
            I => \N__4512\
        );

    \I__1028\ : SRMux
    port map (
            O => \N__4570\,
            I => \N__4512\
        );

    \I__1027\ : SRMux
    port map (
            O => \N__4569\,
            I => \N__4512\
        );

    \I__1026\ : SRMux
    port map (
            O => \N__4568\,
            I => \N__4512\
        );

    \I__1025\ : SRMux
    port map (
            O => \N__4567\,
            I => \N__4512\
        );

    \I__1024\ : SRMux
    port map (
            O => \N__4566\,
            I => \N__4512\
        );

    \I__1023\ : SRMux
    port map (
            O => \N__4565\,
            I => \N__4512\
        );

    \I__1022\ : GlobalMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__1021\ : gio2CtrlBuf
    port map (
            O => \N__4509\,
            I => i_rst_c_g
        );

    \I__1020\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__4500\,
            I => \N__4496\
        );

    \I__1017\ : IoInMux
    port map (
            O => \N__4499\,
            I => \N__4493\
        );

    \I__1016\ : Span4Mux_h
    port map (
            O => \N__4496\,
            I => \N__4490\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4493\,
            I => \N__4487\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__4490\,
            I => i_rx_clk_c
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__4487\,
            I => i_rx_clk_c
        );

    \I__1012\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4478\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4469\
        );

    \I__1008\ : Span4Mux_s2_v
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__4469\,
            I => \rx_sampling_clockZ0\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__4466\,
            I => \rx_sampling_clockZ0\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4455\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4455\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4455\,
            I => \N__4449\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4444\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4444\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4441\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__4449\,
            I => \N__4436\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4436\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4441\,
            I => \rx_sampling_clock_reg1_fastZ0\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__4436\,
            I => \rx_sampling_clock_reg1_fastZ0\
        );

    \I__995\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4423\
        );

    \I__994\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4415\
        );

    \I__993\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4415\
        );

    \I__992\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4415\
        );

    \I__991\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4408\
        );

    \I__990\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4408\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4423\,
            I => \N__4405\
        );

    \I__988\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4402\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4399\
        );

    \I__986\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4396\
        );

    \I__985\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4393\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4408\,
            I => \stateZ0Z_10\
        );

    \I__983\ : Odrv12
    port map (
            O => \N__4405\,
            I => \stateZ0Z_10\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4402\,
            I => \stateZ0Z_10\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__4399\,
            I => \stateZ0Z_10\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4396\,
            I => \stateZ0Z_10\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4393\,
            I => \stateZ0Z_10\
        );

    \I__978\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4375\
        );

    \I__977\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4372\
        );

    \I__976\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4369\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4375\,
            I => \N__4366\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4372\,
            I => \rx_clk_regZ0Z1\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4369\,
            I => \rx_clk_regZ0Z1\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__4366\,
            I => \rx_clk_regZ0Z1\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \N__4355\
        );

    \I__970\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4352\
        );

    \I__969\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4349\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4352\,
            I => \rx_clk_regZ0Z2\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4349\,
            I => \rx_clk_regZ0Z2\
        );

    \I__966\ : IoInMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__964\ : Span4Mux_s3_h
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__4335\,
            I => o_framing_error_c
        );

    \I__962\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4323\
        );

    \I__961\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4323\
        );

    \I__960\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4318\
        );

    \I__959\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4318\
        );

    \I__958\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4315\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4312\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4318\,
            I => \N__4309\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4315\,
            I => \clear_line_statusZ0\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__4312\,
            I => \clear_line_statusZ0\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__4309\,
            I => \clear_line_statusZ0\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__951\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4295\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__4298\,
            I => \N__4292\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4295\,
            I => \N__4288\
        );

    \I__948\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4283\
        );

    \I__947\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4283\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__4288\,
            I => \N__4280\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4283\,
            I => \N__4277\
        );

    \I__944\ : Span4Mux_h
    port map (
            O => \N__4280\,
            I => \N__4274\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__4274\,
            I => i_parity_en_c
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4271\,
            I => i_parity_en_c
        );

    \I__940\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__4254\,
            I => i_stick_parity_en_c
        );

    \I__935\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4247\
        );

    \I__934\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4244\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4247\,
            I => \stick_parity_bitZ0\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4244\,
            I => \stick_parity_bitZ0\
        );

    \I__931\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4234\
        );

    \I__930\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4230\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__4237\,
            I => \N__4227\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4224\
        );

    \I__927\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4221\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4230\,
            I => \N__4218\
        );

    \I__925\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4215\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__4224\,
            I => \N__4210\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4221\,
            I => \N__4210\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4218\,
            I => \rx_dataZ0Z_3\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4215\,
            I => \rx_dataZ0Z_3\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__4210\,
            I => \rx_dataZ0Z_3\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__4203\,
            I => \N__4197\
        );

    \I__918\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4194\
        );

    \I__917\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4191\
        );

    \I__916\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4188\
        );

    \I__915\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4185\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4194\,
            I => \N__4182\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4177\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4177\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4185\,
            I => \rx_dataZ0Z_4\
        );

    \I__910\ : Odrv12
    port map (
            O => \N__4182\,
            I => \rx_dataZ0Z_4\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4177\,
            I => \rx_dataZ0Z_4\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__907\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4159\
        );

    \I__905\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4155\
        );

    \I__904\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4152\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__4159\,
            I => \N__4149\
        );

    \I__902\ : InMux
    port map (
            O => \N__4158\,
            I => \N__4146\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4155\,
            I => \N__4141\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4141\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__4149\,
            I => \rx_dataZ0Z_5\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4146\,
            I => \rx_dataZ0Z_5\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__4141\,
            I => \rx_dataZ0Z_5\
        );

    \I__896\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4130\
        );

    \I__895\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4127\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4130\,
            I => \N__4122\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4127\,
            I => \N__4119\
        );

    \I__892\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4116\
        );

    \I__891\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4113\
        );

    \I__890\ : Span4Mux_h
    port map (
            O => \N__4122\,
            I => \N__4110\
        );

    \I__889\ : Sp12to4
    port map (
            O => \N__4119\,
            I => \N__4105\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4105\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4113\,
            I => \rx_dataZ0Z_2\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__4110\,
            I => \rx_dataZ0Z_2\
        );

    \I__885\ : Odrv12
    port map (
            O => \N__4105\,
            I => \rx_dataZ0Z_2\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__4098\,
            I => \N__4092\
        );

    \I__883\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4088\
        );

    \I__882\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4083\
        );

    \I__881\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4083\
        );

    \I__880\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4078\
        );

    \I__879\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4078\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N__4075\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4083\,
            I => \N_103\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4078\,
            I => \N_103\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__4075\,
            I => \N_103\
        );

    \I__874\ : CEMux
    port map (
            O => \N__4068\,
            I => \N__4065\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__872\ : Span4Mux_h
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__4059\,
            I => \N_103_0\
        );

    \I__870\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4050\
        );

    \I__869\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4050\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4050\,
            I => timeout_counter_2_sqmuxa
        );

    \I__867\ : InMux
    port map (
            O => \N__4047\,
            I => \N__4043\
        );

    \I__866\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4040\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4043\,
            I => \rx_sampling_counterZ0Z_2\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4040\,
            I => \rx_sampling_counterZ0Z_2\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__4035\,
            I => \N__4031\
        );

    \I__862\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4023\
        );

    \I__861\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4023\
        );

    \I__860\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4023\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4023\,
            I => \rx_sampling_counterZ0Z_1\
        );

    \I__858\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4017\,
            I => \rx_sampling_counter_RNO_0Z0Z_3\
        );

    \I__856\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4004\
        );

    \I__855\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4004\
        );

    \I__854\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4004\
        );

    \I__853\ : InMux
    port map (
            O => \N__4011\,
            I => \N__4001\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4004\,
            I => \rx_sampling_counterZ0Z_0\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4001\,
            I => \rx_sampling_counterZ0Z_0\
        );

    \I__850\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3991\
        );

    \I__849\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3988\
        );

    \I__848\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3985\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__3991\,
            I => \rx_sampling_counterZ0Z_3\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__3988\,
            I => \rx_sampling_counterZ0Z_3\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__3985\,
            I => \rx_sampling_counterZ0Z_3\
        );

    \I__844\ : ClkMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__843\ : ClkMux
    port map (
            O => \N__3977\,
            I => \N__3972\
        );

    \I__842\ : GlobalMux
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__841\ : gio2CtrlBuf
    port map (
            O => \N__3969\,
            I => i_rx_clk_c_g
        );

    \I__840\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__3960\,
            I => \N__3957\
        );

    \I__837\ : Span4Mux_v
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__3954\,
            I => i_clear_linestatusreg_c
        );

    \I__835\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__3948\,
            I => \N__3944\
        );

    \I__833\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3941\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__3944\,
            I => \N__3936\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__3941\,
            I => \N__3936\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__3930\,
            I => i_start_rx_c
        );

    \I__827\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__3924\,
            I => \N__3920\
        );

    \I__825\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3917\
        );

    \I__824\ : Span4Mux_v
    port map (
            O => \N__3920\,
            I => \N__3910\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__3917\,
            I => \N__3907\
        );

    \I__822\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3900\
        );

    \I__821\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3900\
        );

    \I__820\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3900\
        );

    \I__819\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3897\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__3910\,
            I => \stateZ0Z_0\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__3907\,
            I => \stateZ0Z_0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__3900\,
            I => \stateZ0Z_0\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__3897\,
            I => \stateZ0Z_0\
        );

    \I__814\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3885\,
            I => \N__3880\
        );

    \I__812\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3877\
        );

    \I__811\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3874\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__3880\,
            I => \timeout_counter_beginZ0\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__3877\,
            I => \timeout_counter_beginZ0\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3874\,
            I => \timeout_counter_beginZ0\
        );

    \I__807\ : CEMux
    port map (
            O => \N__3867\,
            I => \N__3864\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__805\ : Odrv12
    port map (
            O => \N__3861\,
            I => \N_42\
        );

    \I__804\ : IoInMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__3855\,
            I => \N__3851\
        );

    \I__802\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3848\
        );

    \I__801\ : Span4Mux_s1_h
    port map (
            O => \N__3851\,
            I => \N__3845\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__3848\,
            I => \N__3842\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__3845\,
            I => \N__3838\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__3842\,
            I => \N__3835\
        );

    \I__797\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3832\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__3838\,
            I => o_break_interrupt_c
        );

    \I__795\ : Odrv4
    port map (
            O => \N__3835\,
            I => o_break_interrupt_c
        );

    \I__794\ : LocalMux
    port map (
            O => \N__3832\,
            I => o_break_interrupt_c
        );

    \I__793\ : IoInMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__791\ : Odrv12
    port map (
            O => \N__3819\,
            I => o_parity_error_c
        );

    \I__790\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__3810\,
            I => \N__3806\
        );

    \I__787\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3803\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__3806\,
            I => \rx_data_ready_regZ0Z1\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3803\,
            I => \rx_data_ready_regZ0Z1\
        );

    \I__784\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3795\,
            I => \N__3792\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__3789\,
            I => \rx_data_ready_regZ0Z2\
        );

    \I__780\ : IoInMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__778\ : Span12Mux_s3_h
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__777\ : Odrv12
    port map (
            O => \N__3777\,
            I => o_rx_data_ready_c
        );

    \I__776\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3770\
        );

    \I__775\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3767\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3757\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3767\,
            I => \N__3757\
        );

    \I__772\ : InMux
    port map (
            O => \N__3766\,
            I => \N__3754\
        );

    \I__771\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3751\
        );

    \I__770\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3746\
        );

    \I__769\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3746\
        );

    \I__768\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3743\
        );

    \I__767\ : Span4Mux_v
    port map (
            O => \N__3757\,
            I => \N__3734\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3754\,
            I => \N__3734\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3751\,
            I => \N__3734\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3746\,
            I => \N__3734\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3743\,
            I => \N__3731\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__3734\,
            I => \N__3728\
        );

    \I__761\ : Span12Mux_v
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__3728\,
            I => \N__3722\
        );

    \I__759\ : Odrv12
    port map (
            O => \N__3725\,
            I => i_no_of_data_bits_c_0
        );

    \I__758\ : Odrv4
    port map (
            O => \N__3722\,
            I => i_no_of_data_bits_c_0
        );

    \I__757\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3713\
        );

    \I__756\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3707\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N__3702\
        );

    \I__754\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3699\
        );

    \I__753\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3696\
        );

    \I__752\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3693\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3707\,
            I => \N__3690\
        );

    \I__750\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3685\
        );

    \I__749\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3685\
        );

    \I__748\ : Span4Mux_v
    port map (
            O => \N__3702\,
            I => \N__3682\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3699\,
            I => \N__3675\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3696\,
            I => \N__3675\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3693\,
            I => \N__3675\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__3690\,
            I => \stateZ0Z_7\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3685\,
            I => \stateZ0Z_7\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__3682\,
            I => \stateZ0Z_7\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__3675\,
            I => \stateZ0Z_7\
        );

    \I__740\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3662\
        );

    \I__739\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3659\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3662\,
            I => \N__3654\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3659\,
            I => \N__3654\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3654\,
            I => \N_181\
        );

    \I__735\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3645\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__3650\,
            I => \N__3641\
        );

    \I__733\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3638\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__3648\,
            I => \N__3632\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3645\,
            I => \N__3628\
        );

    \I__730\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3623\
        );

    \I__729\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3623\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3638\,
            I => \N__3620\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3637\,
            I => \N__3614\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3636\,
            I => \N__3610\
        );

    \I__725\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3607\
        );

    \I__724\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3604\
        );

    \I__723\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3601\
        );

    \I__722\ : Span4Mux_s1_h
    port map (
            O => \N__3628\,
            I => \N__3594\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3594\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__3620\,
            I => \N__3594\
        );

    \I__719\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3591\
        );

    \I__718\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3580\
        );

    \I__717\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3580\
        );

    \I__716\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3580\
        );

    \I__715\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3580\
        );

    \I__714\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3580\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N__3575\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3604\,
            I => \N__3575\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3601\,
            I => \rx_sampling_clock_regZ0Z1\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__3594\,
            I => \rx_sampling_clock_regZ0Z1\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3591\,
            I => \rx_sampling_clock_regZ0Z1\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3580\,
            I => \rx_sampling_clock_regZ0Z1\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__3575\,
            I => \rx_sampling_clock_regZ0Z1\
        );

    \I__706\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3561\,
            I => \N__3553\
        );

    \I__704\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3544\
        );

    \I__703\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3544\
        );

    \I__702\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3544\
        );

    \I__701\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3544\
        );

    \I__700\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3541\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__3553\,
            I => \stateZ0Z_2\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3544\,
            I => \stateZ0Z_2\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3541\,
            I => \stateZ0Z_2\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__3534\,
            I => \N_380_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__693\ : Odrv12
    port map (
            O => \N__3525\,
            I => \N_161\
        );

    \I__692\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N__3516\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__3516\,
            I => \N__3513\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__3513\,
            I => \N_379\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__3510\,
            I => \N__3507\
        );

    \I__687\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3498\
        );

    \I__686\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3495\
        );

    \I__685\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3488\
        );

    \I__684\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3488\
        );

    \I__683\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3488\
        );

    \I__682\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3483\
        );

    \I__681\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3483\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3498\,
            I => \N__3478\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3495\,
            I => \N__3478\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3488\,
            I => \N_142\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3483\,
            I => \N_142\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3478\,
            I => \N_142\
        );

    \I__675\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3465\,
            I => \N_159\
        );

    \I__672\ : CEMux
    port map (
            O => \N__3462\,
            I => \N__3458\
        );

    \I__671\ : CEMux
    port map (
            O => \N__3461\,
            I => \N__3455\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3458\,
            I => \N__3451\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3447\
        );

    \I__668\ : CEMux
    port map (
            O => \N__3454\,
            I => \N__3444\
        );

    \I__667\ : Span4Mux_h
    port map (
            O => \N__3451\,
            I => \N__3441\
        );

    \I__666\ : CEMux
    port map (
            O => \N__3450\,
            I => \N__3438\
        );

    \I__665\ : Sp12to4
    port map (
            O => \N__3447\,
            I => \N__3431\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3444\,
            I => \N__3431\
        );

    \I__663\ : Sp12to4
    port map (
            O => \N__3441\,
            I => \N__3431\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3438\,
            I => \N_16_i\
        );

    \I__661\ : Odrv12
    port map (
            O => \N__3431\,
            I => \N_16_i\
        );

    \I__660\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3420\
        );

    \I__659\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3417\
        );

    \I__658\ : InMux
    port map (
            O => \N__3424\,
            I => \N__3410\
        );

    \I__657\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3407\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3404\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3417\,
            I => \N__3401\
        );

    \I__654\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3396\
        );

    \I__653\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3396\
        );

    \I__652\ : InMux
    port map (
            O => \N__3414\,
            I => \N__3393\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3413\,
            I => \N__3387\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3410\,
            I => \N__3384\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3407\,
            I => \N__3381\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__3404\,
            I => \N__3378\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__3401\,
            I => \N__3371\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3396\,
            I => \N__3371\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3393\,
            I => \N__3371\
        );

    \I__644\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3364\
        );

    \I__643\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3364\
        );

    \I__642\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3364\
        );

    \I__641\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3361\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__3384\,
            I => \N__3356\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__3381\,
            I => \N__3356\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__3378\,
            I => \rx_sampling_clock_regZ0Z2\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__3371\,
            I => \rx_sampling_clock_regZ0Z2\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3364\,
            I => \rx_sampling_clock_regZ0Z2\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3361\,
            I => \rx_sampling_clock_regZ0Z2\
        );

    \I__634\ : Odrv4
    port map (
            O => \N__3356\,
            I => \rx_sampling_clock_regZ0Z2\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3345\,
            I => \N__3342\
        );

    \I__632\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3335\
        );

    \I__631\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3335\
        );

    \I__630\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3332\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3335\,
            I => \N__3327\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3332\,
            I => \N__3323\
        );

    \I__627\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3318\
        );

    \I__626\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3318\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__3327\,
            I => \N__3315\
        );

    \I__624\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3312\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__3323\,
            I => \N__3309\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3318\,
            I => \N__3306\
        );

    \I__621\ : Span4Mux_s1_h
    port map (
            O => \N__3315\,
            I => \N__3301\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3312\,
            I => \N__3301\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__3309\,
            I => \modem_serial_data_fastZ0\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__3306\,
            I => \modem_serial_data_fastZ0\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__3301\,
            I => \modem_serial_data_fastZ0\
        );

    \I__616\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__614\ : Span4Mux_s3_h
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3285\,
            I => \N_88\
        );

    \I__612\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__3276\,
            I => \N__3272\
        );

    \I__609\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3269\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__3272\,
            I => \rx_sampling_startZ0\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3269\,
            I => \rx_sampling_startZ0\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3264\,
            I => \N_103_cascade_\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__3261\,
            I => \o_timeout5_3_cascade_\
        );

    \I__604\ : IoInMux
    port map (
            O => \N__3258\,
            I => \N__3255\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__602\ : IoSpan4Mux
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__601\ : Span4Mux_s2_h
    port map (
            O => \N__3249\,
            I => \N__3246\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__3246\,
            I => \N__3243\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__3243\,
            I => o_timeout_c
        );

    \I__598\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3233\
        );

    \I__597\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3233\
        );

    \I__596\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3230\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3233\,
            I => \timeout_counterZ0Z_0\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3230\,
            I => \timeout_counterZ0Z_0\
        );

    \I__593\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3218\
        );

    \I__592\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3218\
        );

    \I__591\ : InMux
    port map (
            O => \N__3223\,
            I => \N__3215\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3218\,
            I => \timeout_counterZ0Z_1\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3215\,
            I => \timeout_counterZ0Z_1\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3210\,
            I => \N__3206\
        );

    \I__587\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3202\
        );

    \I__586\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3199\
        );

    \I__585\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3196\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3202\,
            I => \timeout_counterZ0Z_2\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3199\,
            I => \timeout_counterZ0Z_2\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3196\,
            I => \timeout_counterZ0Z_2\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__3189\,
            I => \N__3185\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__3188\,
            I => \N__3182\
        );

    \I__579\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3178\
        );

    \I__578\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3175\
        );

    \I__577\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3172\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3178\,
            I => \timeout_counterZ0Z_3\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3175\,
            I => \timeout_counterZ0Z_3\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3172\,
            I => \timeout_counterZ0Z_3\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__3165\,
            I => \o2_cascade_\
        );

    \I__572\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3159\,
            I => \timeout_counter_RNI09R61Z0Z_5\
        );

    \I__570\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3152\
        );

    \I__569\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3149\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3152\,
            I => \N__3144\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3149\,
            I => \N__3144\
        );

    \I__566\ : Span4Mux_h
    port map (
            O => \N__3144\,
            I => \N__3141\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__3141\,
            I => \N__3138\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__3138\,
            I => i_clear_rxdataready_c
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__562\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3129\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__3126\,
            I => timeout_counter_s_4
        );

    \I__559\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3118\
        );

    \I__558\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3113\
        );

    \I__557\ : InMux
    port map (
            O => \N__3121\,
            I => \N__3113\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3118\,
            I => \N__3110\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3113\,
            I => \timeout_counterZ0Z_4\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__3110\,
            I => \timeout_counterZ0Z_4\
        );

    \I__553\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3096\
        );

    \I__552\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3096\
        );

    \I__551\ : InMux
    port map (
            O => \N__3103\,
            I => \N__3093\
        );

    \I__550\ : InMux
    port map (
            O => \N__3102\,
            I => \N__3088\
        );

    \I__549\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3088\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3096\,
            I => \clearrxdatareadyZ0Z1\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3093\,
            I => \clearrxdatareadyZ0Z1\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3088\,
            I => \clearrxdatareadyZ0Z1\
        );

    \I__545\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3074\
        );

    \I__544\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3074\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3079\,
            I => \N__3070\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3074\,
            I => \N__3065\
        );

    \I__541\ : InMux
    port map (
            O => \N__3073\,
            I => \N__3060\
        );

    \I__540\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3060\
        );

    \I__539\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3055\
        );

    \I__538\ : InMux
    port map (
            O => \N__3068\,
            I => \N__3055\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__3065\,
            I => \N_345_0_i\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3060\,
            I => \N_345_0_i\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3055\,
            I => \N_345_0_i\
        );

    \I__534\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__3042\,
            I => timeout_counter_s_5
        );

    \I__531\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3035\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3038\,
            I => \N__3031\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3035\,
            I => \N__3028\
        );

    \I__528\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3023\
        );

    \I__527\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3023\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__3028\,
            I => \timeout_counterZ0Z_5\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3023\,
            I => \timeout_counterZ0Z_5\
        );

    \I__524\ : CEMux
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3015\,
            I => \N__3011\
        );

    \I__522\ : CEMux
    port map (
            O => \N__3014\,
            I => \N__3008\
        );

    \I__521\ : Sp12to4
    port map (
            O => \N__3011\,
            I => \N__3003\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3008\,
            I => \N__3003\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__3003\,
            I => timeout_countere_0_i
        );

    \I__518\ : InMux
    port map (
            O => \N__3000\,
            I => \bfn_4_9_0_\
        );

    \I__517\ : InMux
    port map (
            O => \N__2997\,
            I => timeout_counter_cry_0
        );

    \I__516\ : InMux
    port map (
            O => \N__2994\,
            I => timeout_counter_cry_1
        );

    \I__515\ : InMux
    port map (
            O => \N__2991\,
            I => timeout_counter_cry_2
        );

    \I__514\ : InMux
    port map (
            O => \N__2988\,
            I => timeout_counter_cry_3
        );

    \I__513\ : InMux
    port map (
            O => \N__2985\,
            I => timeout_counter_cry_4
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__2982\,
            I => \N_92_cascade_\
        );

    \I__511\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2973\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__2978\,
            I => \N__2970\
        );

    \I__509\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2963\
        );

    \I__508\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2963\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2973\,
            I => \N__2960\
        );

    \I__506\ : InMux
    port map (
            O => \N__2970\,
            I => \N__2957\
        );

    \I__505\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2952\
        );

    \I__504\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2952\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N_183\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__2960\,
            I => \N_183\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2957\,
            I => \N_183\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2952\,
            I => \N_183\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__2943\,
            I => \N_147_cascade_\
        );

    \I__498\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2928\
        );

    \I__497\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2928\
        );

    \I__496\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2928\
        );

    \I__495\ : InMux
    port map (
            O => \N__2937\,
            I => \N__2925\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__2936\,
            I => \N__2922\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__2935\,
            I => \N__2919\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2928\,
            I => \N__2913\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2925\,
            I => \N__2910\
        );

    \I__490\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2905\
        );

    \I__489\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2905\
        );

    \I__488\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2902\
        );

    \I__487\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2897\
        );

    \I__486\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2897\
        );

    \I__485\ : Span4Mux_v
    port map (
            O => \N__2913\,
            I => \N__2890\
        );

    \I__484\ : Span4Mux_h
    port map (
            O => \N__2910\,
            I => \N__2890\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2905\,
            I => \N__2890\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2902\,
            I => \stateZ0Z_9\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2897\,
            I => \stateZ0Z_9\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__2890\,
            I => \stateZ0Z_9\
        );

    \I__479\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2878\
        );

    \I__478\ : InMux
    port map (
            O => \N__2882\,
            I => \N__2871\
        );

    \I__477\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2871\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2878\,
            I => \N__2868\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__2877\,
            I => \N__2865\
        );

    \I__474\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2861\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2871\,
            I => \N__2856\
        );

    \I__472\ : Span4Mux_v
    port map (
            O => \N__2868\,
            I => \N__2856\
        );

    \I__471\ : InMux
    port map (
            O => \N__2865\,
            I => \N__2851\
        );

    \I__470\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2851\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N_182\
        );

    \I__468\ : Odrv4
    port map (
            O => \N__2856\,
            I => \N_182\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2851\,
            I => \N_182\
        );

    \I__466\ : InMux
    port map (
            O => \N__2844\,
            I => \N__2835\
        );

    \I__465\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2832\
        );

    \I__464\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2829\
        );

    \I__463\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2819\
        );

    \I__462\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2819\
        );

    \I__461\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2819\
        );

    \I__460\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2816\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2835\,
            I => \N__2809\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2832\,
            I => \N__2809\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2829\,
            I => \N__2809\
        );

    \I__456\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2802\
        );

    \I__455\ : InMux
    port map (
            O => \N__2827\,
            I => \N__2802\
        );

    \I__454\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2802\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2819\,
            I => \N__2797\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2797\
        );

    \I__451\ : Span4Mux_v
    port map (
            O => \N__2809\,
            I => \N__2792\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2802\,
            I => \N__2792\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__2797\,
            I => \modem_serial_data_repZ0Z1\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2792\,
            I => \modem_serial_data_repZ0Z1\
        );

    \I__447\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__2781\,
            I => \N_377\
        );

    \I__444\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2771\
        );

    \I__443\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2766\
        );

    \I__442\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2766\
        );

    \I__441\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2763\
        );

    \I__440\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2760\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2771\,
            I => \N__2755\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2766\,
            I => \N__2755\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2763\,
            I => \rx_sampling_clock_reg2_fastZ0\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2760\,
            I => \rx_sampling_clock_reg2_fastZ0\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__2755\,
            I => \rx_sampling_clock_reg2_fastZ0\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__433\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2740\
        );

    \I__432\ : InMux
    port map (
            O => \N__2744\,
            I => \N__2737\
        );

    \I__431\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2733\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2740\,
            I => \N__2728\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2737\,
            I => \N__2728\
        );

    \I__428\ : InMux
    port map (
            O => \N__2736\,
            I => \N__2722\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2733\,
            I => \N__2719\
        );

    \I__426\ : Span4Mux_v
    port map (
            O => \N__2728\,
            I => \N__2716\
        );

    \I__425\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2711\
        );

    \I__424\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2711\
        );

    \I__423\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2708\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2722\,
            I => \N__2703\
        );

    \I__421\ : Span4Mux_s1_h
    port map (
            O => \N__2719\,
            I => \N__2703\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2716\,
            I => \stateZ0Z_5\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2711\,
            I => \stateZ0Z_5\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2708\,
            I => \stateZ0Z_5\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__2703\,
            I => \stateZ0Z_5\
        );

    \I__416\ : InMux
    port map (
            O => \N__2694\,
            I => \N__2689\
        );

    \I__415\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2686\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2692\,
            I => \N__2682\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2689\,
            I => \N__2675\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2686\,
            I => \N__2675\
        );

    \I__411\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2672\
        );

    \I__410\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2669\
        );

    \I__409\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2666\
        );

    \I__408\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2663\
        );

    \I__407\ : Span4Mux_s1_h
    port map (
            O => \N__2675\,
            I => \N__2660\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2672\,
            I => \stateZ0Z_4\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2669\,
            I => \stateZ0Z_4\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2666\,
            I => \stateZ0Z_4\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2663\,
            I => \stateZ0Z_4\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__2660\,
            I => \stateZ0Z_4\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__2649\,
            I => \N__2646\
        );

    \I__400\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2636\
        );

    \I__399\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2636\
        );

    \I__398\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2631\
        );

    \I__397\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2631\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__2642\,
            I => \N__2628\
        );

    \I__395\ : InMux
    port map (
            O => \N__2641\,
            I => \N__2625\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2620\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2631\,
            I => \N__2620\
        );

    \I__392\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2617\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2625\,
            I => \stateZ0Z_3\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__2620\,
            I => \stateZ0Z_3\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2617\,
            I => \stateZ0Z_3\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2610\,
            I => \N_143_cascade_\
        );

    \I__387\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2604\,
            I => \N__2600\
        );

    \I__385\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2597\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__2600\,
            I => \N__2594\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2597\,
            I => \rx_dataZ0Z_0\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__2594\,
            I => \rx_dataZ0Z_0\
        );

    \I__381\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2586\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2586\,
            I => \N__2583\
        );

    \I__379\ : Odrv4
    port map (
            O => \N__2583\,
            I => \N_115\
        );

    \I__378\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2573\
        );

    \I__377\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2573\
        );

    \I__376\ : InMux
    port map (
            O => \N__2578\,
            I => \N__2566\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2573\,
            I => \N__2563\
        );

    \I__374\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2560\
        );

    \I__373\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2553\
        );

    \I__372\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2553\
        );

    \I__371\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2553\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2566\,
            I => \N_174\
        );

    \I__369\ : Odrv4
    port map (
            O => \N__2563\,
            I => \N_174\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2560\,
            I => \N_174\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2553\,
            I => \N_174\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__2544\,
            I => \N_150_cascade_\
        );

    \I__365\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2538\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2538\,
            I => rx_data_35_0_iv_0_a2_0_1_4
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__2535\,
            I => \N_142_cascade_\
        );

    \I__362\ : InMux
    port map (
            O => \N__2532\,
            I => \N__2529\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2529\,
            I => \N_155\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__2526\,
            I => \rx_data_RNO_2Z0Z_1_cascade_\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2523\,
            I => \rx_data_RNO_1Z0Z_1_cascade_\
        );

    \I__358\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2517\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2517\,
            I => \N__2514\
        );

    \I__356\ : Odrv4
    port map (
            O => \N__2514\,
            I => rx_data_35_0_i_1_1
        );

    \I__355\ : CEMux
    port map (
            O => \N__2511\,
            I => \N__2508\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2508\,
            I => \N__2505\
        );

    \I__353\ : Span4Mux_v
    port map (
            O => \N__2505\,
            I => \N__2502\
        );

    \I__352\ : Odrv4
    port map (
            O => \N__2502\,
            I => un1_framing_error_0_sqmuxa_0_i
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__2499\,
            I => \N_13_i_1_1_cascade_\
        );

    \I__350\ : InMux
    port map (
            O => \N__2496\,
            I => \N__2491\
        );

    \I__349\ : InMux
    port map (
            O => \N__2495\,
            I => \N__2486\
        );

    \I__348\ : InMux
    port map (
            O => \N__2494\,
            I => \N__2486\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2491\,
            I => \N__2483\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2486\,
            I => \clear_data_readyZ0\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__2483\,
            I => \clear_data_readyZ0\
        );

    \I__344\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2475\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2475\,
            I => \N_386\
        );

    \I__342\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2466\
        );

    \I__341\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2466\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2466\,
            I => \N__2463\
        );

    \I__339\ : Odrv4
    port map (
            O => \N__2463\,
            I => \N_13_i_1\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2460\,
            I => \N_165_cascade_\
        );

    \I__337\ : InMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2454\,
            I => rx_data_35_0_iv_0_a2_1_0_0
        );

    \I__335\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2448\,
            I => break_interrupt_e_sn
        );

    \I__333\ : InMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2442\,
            I => break_interrupt_e_rn_0
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__2439\,
            I => \break_interrupt_0_sqmuxa_0_a2_6_cascade_\
        );

    \I__330\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2433\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2433\,
            I => break_interrupt_0_sqmuxa_0_a2_7
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2430\,
            I => \un1_rx_data_0_sqmuxa_2_i_a2_d_0_0_cascade_\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2427\,
            I => \rx_data_35_0_iv_0_a2_0_0_4_cascade_\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2424\,
            I => \N__2418\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2423\,
            I => \N__2415\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2422\,
            I => \N__2412\
        );

    \I__323\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2407\
        );

    \I__322\ : InMux
    port map (
            O => \N__2418\,
            I => \N__2407\
        );

    \I__321\ : InMux
    port map (
            O => \N__2415\,
            I => \N__2401\
        );

    \I__320\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2398\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2407\,
            I => \N__2395\
        );

    \I__318\ : InMux
    port map (
            O => \N__2406\,
            I => \N__2392\
        );

    \I__317\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2387\
        );

    \I__316\ : InMux
    port map (
            O => \N__2404\,
            I => \N__2387\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2401\,
            I => \N__2382\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2398\,
            I => \N__2382\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__2395\,
            I => \N__2375\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2392\,
            I => \N__2375\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2387\,
            I => \N__2375\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__2382\,
            I => \N__2370\
        );

    \I__309\ : Span4Mux_v
    port map (
            O => \N__2375\,
            I => \N__2370\
        );

    \I__308\ : Span4Mux_v
    port map (
            O => \N__2370\,
            I => \N__2367\
        );

    \I__307\ : Odrv4
    port map (
            O => \N__2367\,
            I => i_no_of_data_bits_c_1
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2364\,
            I => \N__2358\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__2363\,
            I => \N__2353\
        );

    \I__304\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2350\
        );

    \I__303\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2347\
        );

    \I__302\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2344\
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__2357\,
            I => \N__2339\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2356\,
            I => \N__2336\
        );

    \I__299\ : InMux
    port map (
            O => \N__2353\,
            I => \N__2333\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2350\,
            I => \N__2330\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2347\,
            I => \N__2325\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2344\,
            I => \N__2325\
        );

    \I__295\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2316\
        );

    \I__294\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2316\
        );

    \I__293\ : InMux
    port map (
            O => \N__2339\,
            I => \N__2316\
        );

    \I__292\ : InMux
    port map (
            O => \N__2336\,
            I => \N__2316\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2333\,
            I => \N__2313\
        );

    \I__290\ : Odrv12
    port map (
            O => \N__2330\,
            I => \stateZ0Z_8\
        );

    \I__289\ : Odrv4
    port map (
            O => \N__2325\,
            I => \stateZ0Z_8\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2316\,
            I => \stateZ0Z_8\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__2313\,
            I => \stateZ0Z_8\
        );

    \I__286\ : CascadeMux
    port map (
            O => \N__2304\,
            I => \N__2299\
        );

    \I__285\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2288\
        );

    \I__284\ : InMux
    port map (
            O => \N__2302\,
            I => \N__2288\
        );

    \I__283\ : InMux
    port map (
            O => \N__2299\,
            I => \N__2288\
        );

    \I__282\ : InMux
    port map (
            O => \N__2298\,
            I => \N__2288\
        );

    \I__281\ : InMux
    port map (
            O => \N__2297\,
            I => \N__2285\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2288\,
            I => \state_fastZ0Z_6\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2285\,
            I => \state_fastZ0Z_6\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2280\,
            I => \N__2276\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2279\,
            I => \N__2273\
        );

    \I__276\ : InMux
    port map (
            O => \N__2276\,
            I => \N__2268\
        );

    \I__275\ : InMux
    port map (
            O => \N__2273\,
            I => \N__2263\
        );

    \I__274\ : InMux
    port map (
            O => \N__2272\,
            I => \N__2263\
        );

    \I__273\ : InMux
    port map (
            O => \N__2271\,
            I => \N__2260\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2268\,
            I => \N__2255\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2263\,
            I => \N__2255\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2260\,
            I => \stateZ0Z_6\
        );

    \I__269\ : Odrv12
    port map (
            O => \N__2255\,
            I => \stateZ0Z_6\
        );

    \I__268\ : InMux
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2247\,
            I => \N__2244\
        );

    \I__266\ : Span4Mux_v
    port map (
            O => \N__2244\,
            I => \N__2241\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2241\,
            I => \N_378\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2238\,
            I => \N__2232\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2237\,
            I => \N__2223\
        );

    \I__262\ : InMux
    port map (
            O => \N__2236\,
            I => \N__2209\
        );

    \I__261\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2209\
        );

    \I__260\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2209\
        );

    \I__259\ : InMux
    port map (
            O => \N__2231\,
            I => \N__2209\
        );

    \I__258\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2209\
        );

    \I__257\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2209\
        );

    \I__256\ : InMux
    port map (
            O => \N__2228\,
            I => \N__2202\
        );

    \I__255\ : InMux
    port map (
            O => \N__2227\,
            I => \N__2202\
        );

    \I__254\ : InMux
    port map (
            O => \N__2226\,
            I => \N__2202\
        );

    \I__253\ : InMux
    port map (
            O => \N__2223\,
            I => \N__2197\
        );

    \I__252\ : InMux
    port map (
            O => \N__2222\,
            I => \N__2197\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2209\,
            I => \N__2190\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2202\,
            I => \N__2190\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2197\,
            I => \N__2190\
        );

    \I__248\ : Span4Mux_v
    port map (
            O => \N__2190\,
            I => \N__2187\
        );

    \I__247\ : Odrv4
    port map (
            O => \N__2187\,
            I => \data_validationZ0\
        );

    \I__246\ : CascadeMux
    port map (
            O => \N__2184\,
            I => \rx_data_35_0_iv_0_a2_0_1_s_0_7_cascade_\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__2181\,
            I => \N_183_cascade_\
        );

    \I__244\ : InMux
    port map (
            O => \N__2178\,
            I => \N__2175\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2175\,
            I => rx_data_35_0_iv_0_a2_0_1_s_0_0_9
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2172\,
            I => \rx_data_35_0_iv_0_a2_0_1_s_0_0_9_cascade_\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__2169\,
            I => \state_ns_i_i_0_a2_0_8_cascade_\
        );

    \I__240\ : InMux
    port map (
            O => \N__2166\,
            I => \N__2163\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2163\,
            I => \N_176\
        );

    \I__238\ : InMux
    port map (
            O => \N__2160\,
            I => \N__2157\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2157\,
            I => rx_data_35_0_iv_0_a2_0_1_3
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__2154\,
            I => \N_148_cascade_\
        );

    \I__235\ : InMux
    port map (
            O => \N__2151\,
            I => \N__2148\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2148\,
            I => rx_data_35_0_iv_0_a2_0_1_5
        );

    \I__233\ : CascadeMux
    port map (
            O => \N__2145\,
            I => \N_152_cascade_\
        );

    \I__232\ : CascadeMux
    port map (
            O => \N__2142\,
            I => \N_157_cascade_\
        );

    \I__231\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2133\
        );

    \I__230\ : InMux
    port map (
            O => \N__2138\,
            I => \N__2133\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2133\,
            I => rx_data_35_0_iv_0_a2_3_out_0
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__2130\,
            I => \N__2127\
        );

    \I__227\ : InMux
    port map (
            O => \N__2127\,
            I => \N__2124\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2124\,
            I => rx_data_35_0_iv_0_a2_0_1_s_0_7
        );

    \I__225\ : InMux
    port map (
            O => \N__2121\,
            I => \N__2116\
        );

    \I__224\ : InMux
    port map (
            O => \N__2120\,
            I => \N__2111\
        );

    \I__223\ : InMux
    port map (
            O => \N__2119\,
            I => \N__2111\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2116\,
            I => i_serial_data_c
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2111\,
            I => i_serial_data_c
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__2106\,
            I => \N__2102\
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__2105\,
            I => \N__2098\
        );

    \I__218\ : InMux
    port map (
            O => \N__2102\,
            I => \N__2091\
        );

    \I__217\ : InMux
    port map (
            O => \N__2101\,
            I => \N__2091\
        );

    \I__216\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2091\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2091\,
            I => i_loopback_en_c
        );

    \I__214\ : InMux
    port map (
            O => \N__2088\,
            I => \N__2083\
        );

    \I__213\ : InMux
    port map (
            O => \N__2087\,
            I => \N__2078\
        );

    \I__212\ : InMux
    port map (
            O => \N__2086\,
            I => \N__2078\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2083\,
            I => i_int_serial_data_c
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2078\,
            I => i_int_serial_data_c
        );

    \I__209\ : CascadeMux
    port map (
            O => \N__2073\,
            I => \N__2070\
        );

    \I__208\ : InMux
    port map (
            O => \N__2070\,
            I => \N__2067\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2067\,
            I => \N__2064\
        );

    \I__206\ : Odrv4
    port map (
            O => \N__2064\,
            I => state_ns_i_i_a2_0_9
        );

    \I__205\ : IoInMux
    port map (
            O => \N__2061\,
            I => \N__2058\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2058\,
            I => \N__2055\
        );

    \I__203\ : Span4Mux_s0_h
    port map (
            O => \N__2055\,
            I => \N__2052\
        );

    \I__202\ : Odrv4
    port map (
            O => \N__2052\,
            I => o_rx_data_c_3
        );

    \I__201\ : IoInMux
    port map (
            O => \N__2049\,
            I => \N__2046\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2046\,
            I => \N__2043\
        );

    \I__199\ : IoSpan4Mux
    port map (
            O => \N__2043\,
            I => \N__2040\
        );

    \I__198\ : Odrv4
    port map (
            O => \N__2040\,
            I => o_rx_data_c_5
        );

    \I__197\ : InMux
    port map (
            O => \N__2037\,
            I => \N__2034\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__2034\,
            I => \N__2031\
        );

    \I__195\ : Odrv4
    port map (
            O => \N__2031\,
            I => \N_187\
        );

    \I__194\ : CascadeMux
    port map (
            O => \N__2028\,
            I => \N_176_cascade_\
        );

    \I__193\ : IoInMux
    port map (
            O => \N__2025\,
            I => \N__2022\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2022\,
            I => o_rx_data_c_6
        );

    \I__191\ : IoInMux
    port map (
            O => \N__2019\,
            I => \N__2016\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__2016\,
            I => o_rx_data_c_7
        );

    \I__189\ : IoInMux
    port map (
            O => \N__2013\,
            I => \N__2010\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__2010\,
            I => \N__2007\
        );

    \I__187\ : Span4Mux_s0_h
    port map (
            O => \N__2007\,
            I => \N__2004\
        );

    \I__186\ : Span4Mux_v
    port map (
            O => \N__2004\,
            I => \N__2001\
        );

    \I__185\ : Odrv4
    port map (
            O => \N__2001\,
            I => o_rx_data_c_1
        );

    \I__184\ : IoInMux
    port map (
            O => \N__1998\,
            I => \N__1995\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1995\,
            I => \N__1992\
        );

    \I__182\ : IoSpan4Mux
    port map (
            O => \N__1992\,
            I => \N__1989\
        );

    \I__181\ : Odrv4
    port map (
            O => \N__1989\,
            I => o_rx_data_c_2
        );

    \I__180\ : IoInMux
    port map (
            O => \N__1986\,
            I => \N__1983\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1983\,
            I => \N__1980\
        );

    \I__178\ : Span4Mux_s0_h
    port map (
            O => \N__1980\,
            I => \N__1977\
        );

    \I__177\ : Span4Mux_v
    port map (
            O => \N__1977\,
            I => \N__1974\
        );

    \I__176\ : Odrv4
    port map (
            O => \N__1974\,
            I => o_rx_data_c_0
        );

    \I__175\ : IoInMux
    port map (
            O => \N__1971\,
            I => \N__1968\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1968\,
            I => \N__1965\
        );

    \I__173\ : IoSpan4Mux
    port map (
            O => \N__1965\,
            I => \N__1962\
        );

    \I__172\ : Odrv4
    port map (
            O => \N__1962\,
            I => o_rx_data_c_4
        );

    \I__171\ : IoInMux
    port map (
            O => \N__1959\,
            I => \N__1956\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1956\,
            I => \N__1953\
        );

    \I__169\ : Span4Mux_s3_h
    port map (
            O => \N__1953\,
            I => \N__1950\
        );

    \I__168\ : Span4Mux_v
    port map (
            O => \N__1950\,
            I => \N__1947\
        );

    \I__167\ : Odrv4
    port map (
            O => \N__1947\,
            I => i_rst_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \i_rst_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1959\,
            GLOBALBUFFEROUTPUT => i_rst_c_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \i_rx_clk_ibuf_RNIGJ1D\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4499\,
            GLOBALBUFFEROUTPUT => i_rx_clk_c_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \state_RNO_0_9_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2405\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3764\,
            lcout => state_ns_i_i_a2_0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_RNO_0_7_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3763\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2404\,
            lcout => \N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_rx_dataZ0Z_6_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2406\,
            in1 => \N__2235\,
            in2 => \_gnd_net_\,
            in3 => \N__4238\,
            lcout => o_rx_data_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \o_rx_dataZ0Z_7_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2236\,
            in1 => \N__3765\,
            in2 => \N__2422\,
            in3 => \N__4133\,
            lcout => o_rx_data_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \o_rx_dataZ0Z_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2230\,
            in2 => \_gnd_net_\,
            in3 => \N__5316\,
            lcout => o_rx_data_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \o_rx_dataZ0Z_2_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2231\,
            lcout => o_rx_data_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \o_rx_dataZ0Z_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2229\,
            in2 => \_gnd_net_\,
            in3 => \N__5244\,
            lcout => o_rx_data_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \o_rx_dataZ0Z_4_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4163\,
            in1 => \_gnd_net_\,
            in2 => \N__2238\,
            in3 => \_gnd_net_\,
            lcout => o_rx_data_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4660\,
            ce => 'H',
            sr => \N__4565\
        );

    \modem_serial_data_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__2119\,
            in1 => \_gnd_net_\,
            in2 => \N__2105\,
            in3 => \N__2086\,
            lcout => \modem_serial_dataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \modem_serial_data_fast_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2121\,
            in1 => \N__2088\,
            in2 => \_gnd_net_\,
            in3 => \N__2101\,
            lcout => \modem_serial_data_fastZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \modem_serial_data_rep1_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__2120\,
            in1 => \_gnd_net_\,
            in2 => \N__2106\,
            in3 => \N__2087\,
            lcout => \modem_serial_data_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \state_9_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__2918\,
            in1 => \N__2362\,
            in2 => \N__2073\,
            in3 => \N__5124\,
            lcout => \stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \o_rx_dataZ0Z_3_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4984\,
            in2 => \_gnd_net_\,
            in3 => \N__2226\,
            lcout => o_rx_data_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \rx_data_ready_reg1_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rx_data_ready_regZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \rx_data_ready_reg2_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3809\,
            lcout => \rx_data_ready_regZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \o_rx_dataZ0Z_5_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__2227\,
            in1 => \N__3766\,
            in2 => \N__2423\,
            in3 => \N__4201\,
            lcout => o_rx_data_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4657\,
            ce => 'H',
            sr => \N__4566\
        );

    \state_7_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__3706\,
            in1 => \N__2037\,
            in2 => \N__2279\,
            in3 => \N__5099\,
            lcout => \stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4659\,
            ce => 'H',
            sr => \N__4567\
        );

    \state_RNIB69F_7_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__4908\,
            in1 => \N__3705\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_176\,
            ltout => \N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_3_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2272\,
            in1 => \N__2917\,
            in2 => \N__2028\,
            in3 => \N__5098\,
            lcout => rx_data_35_0_iv_0_a2_0_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_5_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2916\,
            in1 => \N__5097\,
            in2 => \N__2364\,
            in3 => \N__2166\,
            lcout => rx_data_35_0_iv_0_a2_0_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_0_3_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__2839\,
            in1 => \N__2361\,
            in2 => \N__4237\,
            in3 => \N__5103\,
            lcout => OPEN,
            ltout => \N_148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_3_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__2160\,
            in1 => \N__3503\,
            in2 => \N__2154\,
            in3 => \N__2138\,
            lcout => \rx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4661\,
            ce => \N__3450\,
            sr => \N__4569\
        );

    \rx_data_RNO_0_5_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__2840\,
            in1 => \N__4158\,
            in2 => \N__2280\,
            in3 => \N__5104\,
            lcout => OPEN,
            ltout => \N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_5_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__2151\,
            in1 => \N__3504\,
            in2 => \N__2145\,
            in3 => \N__2139\,
            lcout => \rx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4661\,
            ce => \N__3450\,
            sr => \N__4569\
        );

    \rx_data_RNO_0_7_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2979\,
            in1 => \N__2744\,
            in2 => \N__2130\,
            in3 => \N__2572\,
            lcout => OPEN,
            ltout => \N_157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_7_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__2250\,
            in1 => \N__5268\,
            in2 => \N__2142\,
            in3 => \N__3505\,
            lcout => \rx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4661\,
            ce => \N__3450\,
            sr => \N__4569\
        );

    \state_RNID3IS1_10_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__2841\,
            in1 => \N__2883\,
            in2 => \_gnd_net_\,
            in3 => \N__4422\,
            lcout => rx_data_35_0_iv_0_a2_3_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_3_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__3559\,
            in1 => \N__3426\,
            in2 => \N__2649\,
            in3 => \N__3651\,
            lcout => \stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4664\,
            ce => 'H',
            sr => \N__4571\
        );

    \modem_serial_data_fast_RNIELQ21_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2641\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__3557\,
            lcout => rx_data_35_0_iv_0_a2_0_1_s_0_7,
            ltout => \rx_data_35_0_iv_0_a2_0_1_s_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_0_6_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2694\,
            in1 => \N__2969\,
            in2 => \N__2184\,
            in3 => \N__2571\,
            lcout => \N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_fast_RNIOI531_6_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4904\,
            in1 => \N__3710\,
            in2 => \N__2363\,
            in3 => \N__2297\,
            lcout => \N_183\,
            ltout => \N_183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_0_8_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3558\,
            in1 => \N__2178\,
            in2 => \N__2181\,
            in3 => \N__2570\,
            lcout => \N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \modem_serial_data_fast_RNIIPQ21_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2693\,
            in1 => \N__3330\,
            in2 => \_gnd_net_\,
            in3 => \N__2743\,
            lcout => rx_data_35_0_iv_0_a2_0_1_s_0_0_9,
            ltout => \rx_data_35_0_iv_0_a2_0_1_s_0_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_0_9_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2645\,
            in1 => \N__2968\,
            in2 => \N__2172\,
            in3 => \N__2569\,
            lcout => \N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_2_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__4755\,
            in1 => \N__5117\,
            in2 => \N__4825\,
            in3 => \N__3560\,
            lcout => \stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4664\,
            ce => 'H',
            sr => \N__4571\
        );

    \state_RNO_0_8_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__3773\,
            in1 => \_gnd_net_\,
            in2 => \N__2424\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \state_ns_i_i_0_a2_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_8_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__3712\,
            in1 => \N__5129\,
            in2 => \N__2169\,
            in3 => \N__2343\,
            lcout => \stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4667\,
            ce => 'H',
            sr => \N__4574\
        );

    \rx_data_RNO_2_4_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__4937\,
            in1 => \_gnd_net_\,
            in2 => \N__2357\,
            in3 => \N__2302\,
            lcout => OPEN,
            ltout => \rx_data_35_0_iv_0_a2_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_4_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2844\,
            in2 => \N__2427\,
            in3 => \N__2876\,
            lcout => rx_data_35_0_iv_0_a2_0_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_fast_6_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__3416\,
            in1 => \N__2303\,
            in2 => \N__2748\,
            in3 => \N__3644\,
            lcout => \state_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4667\,
            ce => 'H',
            sr => \N__4574\
        );

    \rx_data_RNO_2_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2342\,
            in2 => \N__2304\,
            in3 => \N__3711\,
            lcout => rx_data_35_0_iv_0_a2_1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_fast_RNIE4LE1_6_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000011011"
        )
    port map (
            in0 => \N__2421\,
            in1 => \N__3774\,
            in2 => \N__2356\,
            in3 => \N__2298\,
            lcout => \N_13_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_6_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__2736\,
            in1 => \N__2271\,
            in2 => \N__3650\,
            in3 => \N__3415\,
            lcout => \stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4667\,
            ce => 'H',
            sr => \N__4574\
        );

    \data_validation_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \data_validationZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4670\,
            ce => \N__2511\,
            sr => \N__4578\
        );

    \rx_data_RNO_1_7_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__3619\,
            in1 => \N__2838\,
            in2 => \N__3413\,
            in3 => \N__2681\,
            lcout => \N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \break_interrupt_RNO_1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4162\,
            in1 => \N__4233\,
            in2 => \N__4986\,
            in3 => \N__4126\,
            lcout => break_interrupt_0_sqmuxa_0_a2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \break_interrupt_RNO_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3841\,
            in1 => \N__2222\,
            in2 => \_gnd_net_\,
            in3 => \N__4329\,
            lcout => break_interrupt_e_rn_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \break_interrupt_RNO_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4330\,
            in1 => \N__2607\,
            in2 => \N__2237\,
            in3 => \N__5200\,
            lcout => break_interrupt_e_sn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \break_interrupt_RNO_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4200\,
            in1 => \N__5315\,
            in2 => \N__5243\,
            in3 => \N__5279\,
            lcout => OPEN,
            ltout => \break_interrupt_0_sqmuxa_0_a2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \break_interrupt_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__2451\,
            in1 => \N__2445\,
            in2 => \N__2439\,
            in3 => \N__2436\,
            lcout => o_break_interrupt_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4658\,
            ce => 'H',
            sr => \N__4568\
        );

    \state_1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__3916\,
            in1 => \N__4793\,
            in2 => \N__4746\,
            in3 => \N__5076\,
            lcout => \stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4662\,
            ce => 'H',
            sr => \N__4570\
        );

    \clear_data_ready_RNI77K81_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__3913\,
            in1 => \N__2494\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => OPEN,
            ltout => \un1_rx_data_0_sqmuxa_2_i_a2_d_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_RNIGRAC2_1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__4727\,
            in1 => \N__4790\,
            in2 => \N__2430\,
            in3 => \N__5072\,
            lcout => \N_16_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clear_data_ready_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__3155\,
            in1 => \N__3947\,
            in2 => \_gnd_net_\,
            in3 => \N__2495\,
            lcout => \clear_data_readyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4662\,
            ce => 'H',
            sr => \N__4570\
        );

    \state_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3425\,
            in1 => \N__3635\,
            in2 => \_gnd_net_\,
            in3 => \N__4925\,
            lcout => \stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4662\,
            ce => 'H',
            sr => \N__4570\
        );

    \timeout_counter_begin_RNO_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__4791\,
            in1 => \N__4728\,
            in2 => \N__5110\,
            in3 => \N__3914\,
            lcout => \N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_start_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__3915\,
            in1 => \N__3275\,
            in2 => \N__4745\,
            in3 => \N__4792\,
            lcout => \rx_sampling_startZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4662\,
            ce => 'H',
            sr => \N__4570\
        );

    \data_validation_RNO_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__4909\,
            in1 => \N__4735\,
            in2 => \N__5113\,
            in3 => \N__2478\,
            lcout => un1_framing_error_0_sqmuxa_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_RNO_0_11_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000110011"
        )
    port map (
            in0 => \N__4426\,
            in1 => \N__4910\,
            in2 => \N__4298\,
            in3 => \N__5086\,
            lcout => OPEN,
            ltout => \N_13_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_11_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__2472\,
            in1 => \N__3666\,
            in2 => \N__2499\,
            in3 => \N__2578\,
            lcout => \stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4665\,
            ce => 'H',
            sr => \N__4572\
        );

    \data_validation_RNO_0_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__2496\,
            in1 => \N__3326\,
            in2 => \N__4926\,
            in3 => \_gnd_net_\,
            lcout => \N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_clock_reg1_fast_RNIL7FA_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__2776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4453\,
            lcout => \N_18_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_RNO_0_10_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__5106\,
            in1 => \N__3665\,
            in2 => \N__2936\,
            in3 => \N__2471\,
            lcout => OPEN,
            ltout => \N_165_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_10_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__5087\,
            in1 => \N__4291\,
            in2 => \N__2460\,
            in3 => \N__4427\,
            lcout => \stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4665\,
            ce => 'H',
            sr => \N__4572\
        );

    \rx_sampling_clock_reg1_fast_RNI1FOP_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4454\,
            in1 => \N__2777\,
            in2 => \N__2935\,
            in3 => \N__4413\,
            lcout => \N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2579\,
            in1 => \N__2828\,
            in2 => \N__2877\,
            in3 => \N__2457\,
            lcout => OPEN,
            ltout => \N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_0_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__3501\,
            in1 => \N__2603\,
            in2 => \N__2610\,
            in3 => \N__2589\,
            lcout => \rx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4668\,
            ce => \N__3454\,
            sr => \N__4575\
        );

    \rx_data_RNO_0_0_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__2826\,
            in2 => \N__3648\,
            in3 => \N__2778\,
            lcout => \N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_0_4_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__2827\,
            in1 => \N__5105\,
            in2 => \N__4203\,
            in3 => \N__3716\,
            lcout => OPEN,
            ltout => \N_150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_4_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__2580\,
            in1 => \N__3502\,
            in2 => \N__2544\,
            in3 => \N__2541\,
            lcout => \rx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4668\,
            ce => \N__3454\,
            sr => \N__4575\
        );

    \state_RNIM5373_10_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4414\,
            in1 => \N__2937\,
            in2 => \N__2978\,
            in3 => \N__2864\,
            lcout => \N_142\,
            ltout => \N_142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_6_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__4971\,
            in1 => \N__2787\,
            in2 => \N__2535\,
            in3 => \N__2532\,
            lcout => \rx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4668\,
            ce => \N__3454\,
            sr => \N__4575\
        );

    \rx_data_RNO_0_1_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__4428\,
            in1 => \N__2843\,
            in2 => \N__5125\,
            in3 => \N__2881\,
            lcout => rx_data_35_0_i_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_2_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4460\,
            in1 => \N__3341\,
            in2 => \N__5204\,
            in3 => \N__4429\,
            lcout => OPEN,
            ltout => \rx_data_RNO_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_1_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5199\,
            in2 => \N__2526\,
            in3 => \N__3414\,
            lcout => OPEN,
            ltout => \rx_data_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__2939\,
            in1 => \N__2977\,
            in2 => \N__2523\,
            in3 => \N__2520\,
            lcout => \rx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4671\,
            ce => \N__3461\,
            sr => \N__4579\
        );

    \rx_data_RNO_2_2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__2775\,
            in1 => \N__4461\,
            in2 => \N__3345\,
            in3 => \N__2938\,
            lcout => OPEN,
            ltout => \N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_2_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2882\,
            in1 => \N__4430\,
            in2 => \N__2982\,
            in3 => \N__2976\,
            lcout => OPEN,
            ltout => \N_147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_2_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__4125\,
            in1 => \N__3294\,
            in2 => \N__2943\,
            in3 => \N__2940\,
            lcout => \rx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4671\,
            ce => \N__3461\,
            sr => \N__4579\
        );

    \state_RNIIBKK1_2_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2725\,
            in1 => \N__2680\,
            in2 => \N__2642\,
            in3 => \N__3556\,
            lcout => \N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_6_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__2842\,
            in1 => \N__2726\,
            in2 => \N__3636\,
            in3 => \N__2774\,
            lcout => \N_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_clock_reg2_fast_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3618\,
            lcout => \rx_sampling_clock_reg2_fastZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4674\,
            ce => 'H',
            sr => \N__4582\
        );

    \state_5_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__3617\,
            in1 => \N__2727\,
            in2 => \N__2692\,
            in3 => \N__3392\,
            lcout => \stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4674\,
            ce => 'H',
            sr => \N__4582\
        );

    \state_4_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__2644\,
            in1 => \N__3391\,
            in2 => \N__3637\,
            in3 => \N__2685\,
            lcout => \stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4674\,
            ce => 'H',
            sr => \N__4582\
        );

    \rx_data_RNO_1_8_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3390\,
            in1 => \N__3613\,
            in2 => \N__4826\,
            in3 => \N__2643\,
            lcout => \N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_clock_reg1_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rx_sampling_clock_regZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4677\,
            ce => 'H',
            sr => \N__4585\
        );

    \rx_sampling_clock_reg2_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => \rx_sampling_clock_regZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4677\,
            ce => 'H',
            sr => \N__4585\
        );

    \timeout_counter_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3080\,
            in1 => \N__3238\,
            in2 => \_gnd_net_\,
            in3 => \N__3000\,
            lcout => \timeout_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => timeout_counter_cry_0,
            clk => \N__4663\,
            ce => \N__3018\,
            sr => \N__4573\
        );

    \timeout_counter_1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3068\,
            in1 => \N__3223\,
            in2 => \_gnd_net_\,
            in3 => \N__2997\,
            lcout => \timeout_counterZ0Z_1\,
            ltout => OPEN,
            carryin => timeout_counter_cry_0,
            carryout => timeout_counter_cry_1,
            clk => \N__4663\,
            ce => \N__3018\,
            sr => \N__4573\
        );

    \timeout_counter_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3081\,
            in1 => \N__3205\,
            in2 => \_gnd_net_\,
            in3 => \N__2994\,
            lcout => \timeout_counterZ0Z_2\,
            ltout => OPEN,
            carryin => timeout_counter_cry_1,
            carryout => timeout_counter_cry_2,
            clk => \N__4663\,
            ce => \N__3018\,
            sr => \N__4573\
        );

    \timeout_counter_3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__3069\,
            in1 => \_gnd_net_\,
            in2 => \N__3188\,
            in3 => \N__2991\,
            lcout => \timeout_counterZ0Z_3\,
            ltout => OPEN,
            carryin => timeout_counter_cry_2,
            carryout => timeout_counter_cry_3,
            clk => \N__4663\,
            ce => \N__3018\,
            sr => \N__4573\
        );

    \timeout_counter_RNO_0_4_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3123\,
            in2 => \_gnd_net_\,
            in3 => \N__2988\,
            lcout => timeout_counter_s_4,
            ltout => OPEN,
            carryin => timeout_counter_cry_3,
            carryout => timeout_counter_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \timeout_counter_RNO_0_5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3039\,
            in2 => \_gnd_net_\,
            in3 => \N__2985\,
            lcout => timeout_counter_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_timeout_RNO_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3034\,
            in1 => \N__3122\,
            in2 => \N__3189\,
            in3 => \N__3209\,
            lcout => OPEN,
            ltout => \o_timeout5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_timeoutZ0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__3225\,
            in1 => \N__3240\,
            in2 => \N__3261\,
            in3 => \_gnd_net_\,
            lcout => o_timeout_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4669\,
            ce => 'H',
            sr => \N__4576\
        );

    \timeout_counter_RNIUV411_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3239\,
            in1 => \N__3224\,
            in2 => \N__3210\,
            in3 => \N__3181\,
            lcout => OPEN,
            ltout => \o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \timeout_counter_begin_RNIPR8U2_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100001011"
        )
    port map (
            in0 => \N__3102\,
            in1 => \N__3884\,
            in2 => \N__3165\,
            in3 => \N__3162\,
            lcout => \N_345_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \timeout_counter_RNI09R61_5_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__3103\,
            in1 => \N__3121\,
            in2 => \N__3038\,
            in3 => \N__3883\,
            lcout => \timeout_counter_RNI09R61Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clearrxdataready1_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3156\,
            lcout => \clearrxdatareadyZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4669\,
            ce => 'H',
            sr => \N__4576\
        );

    \rx_clk_reg2_RNIK6ND_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__4358\,
            in1 => \N__4378\,
            in2 => \_gnd_net_\,
            in3 => \N__3101\,
            lcout => timeout_countere_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \timeout_counter_4_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__4055\,
            in1 => \N__3105\,
            in2 => \N__3135\,
            in3 => \N__3073\,
            lcout => \timeout_counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4672\,
            ce => \N__3014\,
            sr => \N__4580\
        );

    \timeout_counter_5_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__3104\,
            in1 => \N__4056\,
            in2 => \N__3079\,
            in3 => \N__3048\,
            lcout => \timeout_counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4672\,
            ce => \N__3014\,
            sr => \N__4580\
        );

    \o_parity_error_obuf_RNO_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3854\,
            lcout => o_parity_error_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_rx_data_ready_obuf_RNO_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3798\,
            lcout => o_rx_data_ready_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_RNI0IHQ_7_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3762\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3717\,
            lcout => \N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_RNO_1_9_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3424\,
            in1 => \N__3649\,
            in2 => \N__4836\,
            in3 => \N__3564\,
            lcout => OPEN,
            ltout => \N_380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_data_9_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__3506\,
            in1 => \N__5229\,
            in2 => \N__3534\,
            in3 => \N__3531\,
            lcout => \rx_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4675\,
            ce => \N__3462\,
            sr => \N__4583\
        );

    \rx_data_8_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__3522\,
            in1 => \N__5308\,
            in2 => \N__3510\,
            in3 => \N__3471\,
            lcout => \rx_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4675\,
            ce => \N__3462\,
            sr => \N__4583\
        );

    \rx_data_RNO_0_2_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__3423\,
            in1 => \N__3340\,
            in2 => \_gnd_net_\,
            in3 => \N__4452\,
            lcout => \N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_start_RNIQR6E_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3927\,
            lcout => \N_103\,
            ltout => \N_103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_counter_RNO_0_3_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__3994\,
            in1 => \N__4046\,
            in2 => \N__3264\,
            in3 => \N__4011\,
            lcout => \rx_sampling_counter_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_clk_reg2_RNID25G_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__4380\,
            in1 => \_gnd_net_\,
            in2 => \N__4359\,
            in3 => \N__3888\,
            lcout => timeout_counter_2_sqmuxa,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_counter_2_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__4014\,
            in1 => \N__4096\,
            in2 => \N__4035\,
            in3 => \N__4047\,
            lcout => \rx_sampling_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3977\,
            ce => 'H',
            sr => \N__4586\
        );

    \rx_sampling_counter_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4030\,
            in2 => \_gnd_net_\,
            in3 => \N__4013\,
            lcout => \rx_sampling_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3977\,
            ce => 'H',
            sr => \N__4586\
        );

    \rx_sampling_counter_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__4034\,
            in1 => \N__3995\,
            in2 => \N__4098\,
            in3 => \N__4020\,
            lcout => \rx_sampling_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3977\,
            ce => 'H',
            sr => \N__4586\
        );

    \rx_sampling_counter_0_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4091\,
            in2 => \_gnd_net_\,
            in3 => \N__4012\,
            lcout => \rx_sampling_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3977\,
            ce => 'H',
            sr => \N__4586\
        );

    \rx_sampling_clock_er_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3996\,
            lcout => \rx_sampling_clockZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3978\,
            ce => \N__4068\,
            sr => \N__4588\
        );

    \clear_line_status_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__3966\,
            in1 => \N__3951\,
            in2 => \_gnd_net_\,
            in3 => \N__4328\,
            lcout => \clear_line_statusZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4666\,
            ce => 'H',
            sr => \N__4577\
        );

    \timeout_counter_begin_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3923\,
            lcout => \timeout_counter_beginZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4673\,
            ce => \N__3867\,
            sr => \N__4581\
        );

    \rx_clk_reg1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rx_clk_regZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4676\,
            ce => 'H',
            sr => \N__4584\
        );

    \rx_sampling_clock_reg1_fast_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4481\,
            lcout => \rx_sampling_clock_reg1_fastZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4676\,
            ce => 'H',
            sr => \N__4584\
        );

    \stick_parity_bit_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__4251\,
            in1 => \N__4431\,
            in2 => \N__4845\,
            in3 => \N__5112\,
            lcout => \stick_parity_bitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4676\,
            ce => 'H',
            sr => \N__4584\
        );

    \rx_clk_reg2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4379\,
            lcout => \rx_clk_regZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4676\,
            ce => 'H',
            sr => \N__4584\
        );

    \o_framing_error_obuf_RNO_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4332\,
            lcout => o_framing_error_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \parity_error_RNO_1_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__4331\,
            in2 => \N__4302\,
            in3 => \N__4939\,
            lcout => parity_error_e_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \parity_error_RNO_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4266\,
            in1 => \N__4250\,
            in2 => \_gnd_net_\,
            in3 => \N__4851\,
            lcout => \N_398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \check_bit_RNO_1_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__4239\,
            in1 => \N__4202\,
            in2 => \N__4170\,
            in3 => \N__4134\,
            lcout => check_bit_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_sampling_clock_sbtinv_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4097\,
            lcout => \N_103_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \check_bit_RNO_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__5301\,
            in1 => \N__5278\,
            in2 => \N__5230\,
            in3 => \N__5205\,
            lcout => check_bit_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \parity_error_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010001001100"
        )
    port map (
            in0 => \N__4946\,
            in1 => \N__5172\,
            in2 => \N__5166\,
            in3 => \N__5154\,
            lcout => \parity_errorZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4679\,
            ce => 'H',
            sr => \N__4589\
        );

    \framing_error_RNO_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__4754\,
            in1 => \N__4927\,
            in2 => \N__4844\,
            in3 => \N__5111\,
            lcout => un1_rx_data_0_sqmuxa_1_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \check_bit_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \N__4992\,
            in2 => \N__4985\,
            in3 => \N__4947\,
            lcout => \check_bitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4680\,
            ce => 'H',
            sr => \N__4590\
        );

    \framing_error_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4843\,
            in2 => \_gnd_net_\,
            in3 => \N__4750\,
            lcout => \framing_errorZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4678\,
            ce => \N__4602\,
            sr => \N__4587\
        );
end \INTERFACE\;
