// ******************************************************************************

// iCEcube Netlister

// Version:            2016.12.27910

// Build Date:         Dec 21 2016 18:07:04

// File Generated:     Mar 12 2017 13:18:20

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "uart" view "INTERFACE"

module uart (
    led,
    test3,
    to_ir,
    test2,
    sd,
    i_serial_data,
    test1,
    o_serial_data,
    from_ir,
    clk_in);

    output [7:0] led;
    output test3;
    output to_ir;
    output test2;
    output sd;
    input i_serial_data;
    output test1;
    output o_serial_data;
    input from_ir;
    input clk_in;

    wire N__6238;
    wire N__6237;
    wire N__6236;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6218;
    wire N__6217;
    wire N__6216;
    wire N__6209;
    wire N__6208;
    wire N__6207;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6191;
    wire N__6190;
    wire N__6189;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6155;
    wire N__6154;
    wire N__6153;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6119;
    wire N__6118;
    wire N__6117;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6101;
    wire N__6100;
    wire N__6099;
    wire N__6092;
    wire N__6091;
    wire N__6090;
    wire N__6073;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6048;
    wire N__6047;
    wire N__6046;
    wire N__6045;
    wire N__6044;
    wire N__6043;
    wire N__6042;
    wire N__6041;
    wire N__6040;
    wire N__6039;
    wire N__6038;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6031;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6022;
    wire N__6021;
    wire N__6020;
    wire N__6019;
    wire N__6018;
    wire N__6017;
    wire N__6016;
    wire N__6015;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5935;
    wire N__5934;
    wire N__5933;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5900;
    wire N__5897;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5599;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5509;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5479;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5451;
    wire N__5448;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5434;
    wire N__5431;
    wire N__5422;
    wire N__5419;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5414;
    wire N__5413;
    wire N__5410;
    wire N__5403;
    wire N__5402;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5377;
    wire N__5368;
    wire N__5367;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5344;
    wire N__5343;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5319;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5287;
    wire N__5284;
    wire N__5279;
    wire N__5272;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5262;
    wire N__5261;
    wire N__5256;
    wire N__5253;
    wire N__5252;
    wire N__5251;
    wire N__5250;
    wire N__5247;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5229;
    wire N__5218;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5191;
    wire N__5190;
    wire N__5189;
    wire N__5188;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5128;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5082;
    wire N__5081;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5042;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5020;
    wire N__5019;
    wire N__5018;
    wire N__5017;
    wire N__5016;
    wire N__5011;
    wire N__5008;
    wire N__5007;
    wire N__5004;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4972;
    wire N__4971;
    wire N__4970;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4951;
    wire N__4948;
    wire N__4939;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4886;
    wire N__4883;
    wire N__4878;
    wire N__4873;
    wire N__4872;
    wire N__4869;
    wire N__4868;
    wire N__4865;
    wire N__4864;
    wire N__4861;
    wire N__4856;
    wire N__4853;
    wire N__4846;
    wire N__4845;
    wire N__4844;
    wire N__4843;
    wire N__4842;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4821;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4777;
    wire N__4774;
    wire N__4773;
    wire N__4772;
    wire N__4771;
    wire N__4766;
    wire N__4761;
    wire N__4756;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4742;
    wire N__4735;
    wire N__4734;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4642;
    wire N__4641;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4626;
    wire N__4623;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4592;
    wire N__4589;
    wire N__4584;
    wire N__4581;
    wire N__4576;
    wire N__4575;
    wire N__4574;
    wire N__4571;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4555;
    wire N__4546;
    wire N__4545;
    wire N__4542;
    wire N__4541;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4525;
    wire N__4516;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4462;
    wire N__4459;
    wire N__4452;
    wire N__4447;
    wire N__4444;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4438;
    wire N__4433;
    wire N__4430;
    wire N__4423;
    wire N__4422;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4393;
    wire N__4386;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4354;
    wire N__4353;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4347;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4315;
    wire N__4314;
    wire N__4309;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4303;
    wire N__4302;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4249;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4245;
    wire N__4244;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4227;
    wire N__4224;
    wire N__4217;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4203;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4195;
    wire N__4190;
    wire N__4189;
    wire N__4188;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4172;
    wire N__4165;
    wire N__4164;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4158;
    wire N__4153;
    wire N__4148;
    wire N__4141;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4100;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4077;
    wire N__4076;
    wire N__4071;
    wire N__4068;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4054;
    wire N__4047;
    wire N__4044;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3994;
    wire N__3991;
    wire N__3990;
    wire N__3989;
    wire N__3988;
    wire N__3983;
    wire N__3978;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3963;
    wire N__3962;
    wire N__3959;
    wire N__3954;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3931;
    wire N__3930;
    wire N__3929;
    wire N__3928;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3916;
    wire N__3913;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3897;
    wire N__3894;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3874;
    wire N__3873;
    wire N__3872;
    wire N__3871;
    wire N__3870;
    wire N__3869;
    wire N__3868;
    wire N__3867;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3840;
    wire N__3839;
    wire N__3838;
    wire N__3837;
    wire N__3834;
    wire N__3825;
    wire N__3822;
    wire N__3817;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3769;
    wire N__3768;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3724;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3712;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3665;
    wire N__3662;
    wire N__3657;
    wire N__3654;
    wire N__3649;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3627;
    wire N__3626;
    wire N__3625;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3609;
    wire N__3608;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3565;
    wire N__3564;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3547;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3535;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3520;
    wire N__3517;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3502;
    wire N__3499;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3484;
    wire N__3481;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3469;
    wire N__3466;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3451;
    wire N__3448;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3433;
    wire N__3430;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3411;
    wire N__3408;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3322;
    wire N__3319;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3283;
    wire N__3280;
    wire N__3279;
    wire N__3274;
    wire N__3271;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3217;
    wire N__3216;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3183;
    wire N__3178;
    wire N__3175;
    wire N__3174;
    wire N__3169;
    wire N__3166;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3148;
    wire N__3147;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3126;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3111;
    wire N__3106;
    wire N__3103;
    wire N__3102;
    wire N__3099;
    wire N__3094;
    wire N__3091;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3079;
    wire N__3078;
    wire N__3073;
    wire N__3070;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3058;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3021;
    wire N__3016;
    wire N__3013;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3001;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2986;
    wire N__2985;
    wire N__2980;
    wire N__2977;
    wire N__2976;
    wire N__2971;
    wire N__2968;
    wire N__2967;
    wire N__2962;
    wire N__2959;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2899;
    wire N__2898;
    wire N__2893;
    wire N__2890;
    wire N__2889;
    wire N__2884;
    wire N__2881;
    wire N__2880;
    wire N__2875;
    wire N__2872;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2854;
    wire N__2853;
    wire N__2848;
    wire N__2845;
    wire N__2844;
    wire N__2839;
    wire N__2836;
    wire N__2835;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2808;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2727;
    wire N__2722;
    wire N__2719;
    wire N__2718;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire \ice_pll_inst.CLKOP ;
    wire GNDG0;
    wire test1_c;
    wire VCCG0;
    wire rst_count_i_19;
    wire o_rx_data_i_6;
    wire shift_reg2Z0Z_14;
    wire shift_reg2Z0Z_13;
    wire shift_reg2Z0Z_15;
    wire shift_reg2Z0Z_11;
    wire shift_reg2Z0Z_10;
    wire shift_reg2Z0Z_12;
    wire shift_reg2Z0Z_9;
    wire shift_reg1Z0Z_1;
    wire shift_reg1Z0Z_2;
    wire rx_rdy_14;
    wire rx_rdy_16_cascade_;
    wire rx_rdy_10;
    wire shift_reg1Z0Z_0;
    wire rx_rdy_11;
    wire shift_reg2Z0Z_4;
    wire shift_reg2Z0Z_5;
    wire shift_reg2Z0Z_6;
    wire shift_reg2Z0Z_7;
    wire shift_reg2Z0Z_8;
    wire GB_BUFFER_clk_in_c_g_THRU_CO;
    wire shift_reg2Z0Z_19;
    wire GB_BUFFER_rst_count_i_g_19_THRU_CO;
    wire shift_reg1Z0Z_8;
    wire shift_reg1Z0Z_9;
    wire shift_reg1Z0Z_15;
    wire shift_reg1Z0Z_10;
    wire shift_reg1Z0Z_14;
    wire shift_reg1Z0Z_13;
    wire shift_reg1Z0Z_11;
    wire shift_reg1Z0Z_12;
    wire shift_reg1Z0Z_7;
    wire i_start_tx_11;
    wire i_start_tx_9;
    wire i_start_tx_8_cascade_;
    wire i_start_tx_10;
    wire shift_reg1Z0Z_5;
    wire shift_reg1Z0Z_6;
    wire shift_reg1Z0Z_3;
    wire shift_reg1Z0Z_4;
    wire un1_rst_countlt18_0;
    wire un1_rst_countlt21_0_i;
    wire shift_reg2Z0Z_17;
    wire shift_reg2Z0Z_16;
    wire shift_reg2Z0Z_18;
    wire shift_reg2Z0Z_0;
    wire rx_rdy_13;
    wire rx_rdy_5;
    wire shift_reg2Z0Z_1;
    wire shift_reg2Z0Z_2;
    wire shift_reg2Z0Z_3;
    wire un1_rst_countlt14_0_cascade_;
    wire un1_rst_countlt17;
    wire bfn_6_3_0_;
    wire rst_countZ0Z_2;
    wire rst_count_1_cry_1;
    wire rst_countZ0Z_3;
    wire rst_count_1_cry_2;
    wire rst_countZ0Z_4;
    wire rst_count_1_cry_3;
    wire rst_countZ0Z_5;
    wire rst_count_1_cry_4;
    wire rst_countZ0Z_6;
    wire rst_count_1_cry_5;
    wire rst_count_1_cry_6;
    wire rst_count_1_cry_7;
    wire rst_count_1_cry_8;
    wire rst_countZ0Z_9;
    wire bfn_6_4_0_;
    wire rst_countZ0Z_10;
    wire rst_count_1_cry_9;
    wire rst_countZ0Z_11;
    wire rst_count_1_cry_10;
    wire rst_countZ0Z_12;
    wire rst_count_1_cry_11;
    wire rst_countZ0Z_13;
    wire rst_count_1_cry_12;
    wire rst_countZ0Z_14;
    wire rst_count_1_cry_13;
    wire rst_countZ0Z_15;
    wire rst_count_1_cry_14;
    wire rst_countZ0Z_16;
    wire rst_count_1_cry_15;
    wire rst_count_1_cry_16;
    wire rst_countZ0Z_17;
    wire bfn_6_5_0_;
    wire rst_countZ0Z_18;
    wire rst_count_1_cry_17;
    wire rst_countZ0Z_19;
    wire rst_count_1_cry_18;
    wire rst_count_1_cry_19;
    wire rst_countZ0Z_20;
    wire rst_countZ0Z_0;
    wire rst_countZ0Z_1;
    wire clk_in_c_g;
    wire un1_rst_countlt21_0_i_g;
    wire o_rx_data_i_5;
    wire bfn_7_1_0_;
    wire un5_count_ext_cry_1;
    wire un5_count_ext_cry_2;
    wire un5_count_ext_cry_3;
    wire count_extZ0Z_3;
    wire count_extZ0Z_1;
    wire count_extZ0Z_2;
    wire from_ir_regZ0Z2;
    wire from_ir_regZ0Z1;
    wire rst_countZ0Z_8;
    wire rst_countZ0Z_7;
    wire un1_rst_countlt9_0;
    wire CONSTANT_ONE_NET;
    wire \uut1.rx_data_35_0_0_6_cascade_ ;
    wire \uut1.N_218_0_cascade_ ;
    wire \uut1.N_217_0_4_cascade_ ;
    wire \uut1.N_216_0_cascade_ ;
    wire count_ext_RNIEM1QZ0Z_1;
    wire count_ext13;
    wire count_extZ0Z_0;
    wire N_95_g;
    wire CLKOS_RNI7KOJZ0Z1;
    wire test2_c;
    wire count_extZ0Z_4;
    wire \uut1.rx_sampling_clock_cnv_1_cascade_ ;
    wire clk_count_RNO_0Z0Z_1_cascade_;
    wire countZ0Z_2;
    wire CLKOS3_3_cascade_;
    wire countZ0Z_1;
    wire countZ0Z_0;
    wire G_7_a0_1;
    wire count_i_3;
    wire CLKOS_i;
    wire G_7_a0_0;
    wire clk_countZ0Z_1;
    wire bfn_8_4_0_;
    wire un3_clk_count_cry_1;
    wire un3_clk_count_cry_2;
    wire un3_clk_count_cry_3;
    wire un3_clk_count_cry_4;
    wire clk_countZ0Z_5;
    wire clk_countZ0Z_2;
    wire clk_count_RNO_0Z0Z_3;
    wire clk_countZ0Z_4;
    wire CLKOS3_3;
    wire clk_countZ0Z_3;
    wire \uut1.rx_data_16_m_6 ;
    wire \uut1.rx_data_13_m_7 ;
    wire \uut1.stateZ0Z_5 ;
    wire \uut1.N_221_0_2_cascade_ ;
    wire \uut1.N_219_0 ;
    wire \uut1.rx_data_22_m_4 ;
    wire \uut1.N_221_0_5_cascade_ ;
    wire \uut1.N_221_0_5 ;
    wire \uut1.stateZ0Z_4 ;
    wire \uut1.N_221_0_2 ;
    wire \uut1.stateZ0Z_6 ;
    wire \uut1.rx_data_25_m_3 ;
    wire \uut1.N_215_0 ;
    wire \uut1.rx_data_19_m_5 ;
    wire \uut1.rx_dataZ0Z_3 ;
    wire \uut1.stateZ0Z_8 ;
    wire \uut1.stateZ0Z_7 ;
    wire \uut1.N_217_0_4 ;
    wire \uut1.N_217_0 ;
    wire \uut1.rx_sampling_clock_RNOZ0 ;
    wire \uut1.CO2 ;
    wire \uut1.N_5 ;
    wire \uut1.rx_sampling_counterZ0Z_2 ;
    wire \uut1.rx_sampling_counterZ0Z_1 ;
    wire \uut1.rx_sampling_counterZ0Z_3 ;
    wire \uut1.rx_sampling_counterZ0Z_0 ;
    wire \uut1.rx_sampling_counter16_cascade_ ;
    wire \uut1.rx_sampling_counter_1_sqmuxa ;
    wire clk_countZ0Z_0;
    wire \uut1.rx_sampling_startZ0 ;
    wire \uut1.rx_data_ready_regZ0Z1 ;
    wire \uut1.rx_data_ready_regZ0Z2 ;
    wire \uut1.rx_dataZ0Z_7 ;
    wire \uut1.state_ns_a2_0_0_2 ;
    wire \uut1.rx_dataZ0Z_6 ;
    wire \uut1.stateZ0Z_1 ;
    wire \uut1.stateZ0Z_11 ;
    wire \uut1.stateZ0Z_0 ;
    wire \uut1.rx_sample_en_cascade_ ;
    wire \uut1.stateZ0Z_3 ;
    wire \uut1.rx_data_10_m_8_cascade_ ;
    wire \uut1.N_220_0 ;
    wire \uut1.rx_dataZ0Z_8 ;
    wire \uut1.rx_sampling_clock_regZ0Z2 ;
    wire \uut1.state_RNID38FZ0Z_1 ;
    wire \uut1.N_221_0 ;
    wire \uut1.rx_dataZ0Z_5 ;
    wire \uut1.rx_sampling_clockZ0 ;
    wire \uut1.rx_sampling_clock_regZ0Z1 ;
    wire \uut1.data_validationZ0 ;
    wire \uut1.rx_dataZ0Z_4 ;
    wire \uut1.modem_serial_dataZ0 ;
    wire \uut1.rx_sample_en ;
    wire \uut1.rx_dataZ0Z_9 ;
    wire \uut1.stateZ0Z_2 ;
    wire \uut1.rx_data_7_m_9 ;
    wire \uut2.stateZ0Z_11 ;
    wire count_RNIH42R1Z0Z_2;
    wire i_start_tx_0;
    wire \uut2.stateZ0Z_0 ;
    wire o_serial_data_c;
    wire \uut2.serial_data_RNOZ0Z_0 ;
    wire \uut2.serial_data_24_iv_3 ;
    wire o_rx_data_6;
    wire \uut2.tx_dataZ0Z_6 ;
    wire \uut2.stateZ0Z_10 ;
    wire \uut2.stateZ0Z_2 ;
    wire \uut2.stateZ0Z_1 ;
    wire \uut2.serial_data_24_iv_2 ;
    wire \uut2.stateZ0Z_13 ;
    wire \uut2.stateZ0Z_3 ;
    wire \uut2.serial_data_24_iv_1 ;
    wire \uut2.stateZ0Z_4 ;
    wire \uut2.serial_data_24_iv_4 ;
    wire o_rx_data_5;
    wire \uut2.tx_dataZ0Z_5 ;
    wire \uut2.tx_dataZ0Z_1 ;
    wire \uut2.tx_dataZ0Z_0 ;
    wire \uut2.tx_dataZ0Z_3 ;
    wire \uut2.stateZ0Z_8 ;
    wire \uut2.stateZ0Z_7 ;
    wire \uut2.tx_dataZ0Z_2 ;
    wire \uut2.stateZ0Z_5 ;
    wire \uut2.stateZ0Z_6 ;
    wire \uut2.tx_dataZ0Z_4 ;
    wire CLKOP_g;
    wire N_123_g;
    wire rst_count_i_g_19;
    wire o_rx_data_3;
    wire o_rx_data_i_3;
    wire o_rx_data_4;
    wire o_rx_data_i_4;
    wire o_rx_data_1;
    wire o_rx_data_i_1;
    wire o_rx_data_2;
    wire o_rx_data_i_2;
    wire o_rx_data_0;
    wire o_rx_data_i_0;
    wire _gnd_net_;

    defparam \ice_pll_inst.ice_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \ice_pll_inst.ice_pll_inst .TEST_MODE=1'b0;
    defparam \ice_pll_inst.ice_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \ice_pll_inst.ice_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \ice_pll_inst.ice_pll_inst .FILTER_RANGE=3'b001;
    defparam \ice_pll_inst.ice_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \ice_pll_inst.ice_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \ice_pll_inst.ice_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \ice_pll_inst.ice_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \ice_pll_inst.ice_pll_inst .DIVR=4'b0000;
    defparam \ice_pll_inst.ice_pll_inst .DIVQ=3'b100;
    defparam \ice_pll_inst.ice_pll_inst .DIVF=7'b0110010;
    defparam \ice_pll_inst.ice_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \ice_pll_inst.ice_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\ice_pll_inst.CLKOP ),
            .REFERENCECLK(N__2941),
            .RESETB(N__3690),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF clk_in_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6236),
            .GLOBALBUFFEROUTPUT(clk_in_c_g));
    IO_PAD clk_in_ibuf_gb_io_iopad (
            .OE(N__6238),
            .DIN(N__6237),
            .DOUT(N__6236),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_gb_io_preio (
            .PADOEN(N__6238),
            .PADOUT(N__6237),
            .PADIN(N__6236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__6227),
            .DIN(N__6226),
            .DOUT(N__6225),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__6227),
            .PADOUT(N__6226),
            .PADIN(N__6225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test1_obuf_iopad (
            .OE(N__6218),
            .DIN(N__6217),
            .DOUT(N__6216),
            .PACKAGEPIN(test1));
    defparam test1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test1_obuf_preio (
            .PADOEN(N__6218),
            .PADOUT(N__6217),
            .PADIN(N__6216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2779),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__6209),
            .DIN(N__6208),
            .DOUT(N__6207),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__6209),
            .PADOUT(N__6208),
            .PADIN(N__6207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5722),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_7_iopad (
            .OE(N__6200),
            .DIN(N__6199),
            .DOUT(N__6198),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__6200),
            .PADOUT(N__6199),
            .PADIN(N__6198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3694),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_4_iopad (
            .OE(N__6191),
            .DIN(N__6190),
            .DOUT(N__6189),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__6191),
            .PADOUT(N__6190),
            .PADIN(N__6189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5791),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test3_obuf_iopad (
            .OE(N__6182),
            .DIN(N__6181),
            .DOUT(N__6180),
            .PACKAGEPIN(test3));
    defparam test3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test3_obuf_preio (
            .PADOEN(N__6182),
            .PADOUT(N__6181),
            .PADIN(N__6180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2920),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__6173),
            .DIN(N__6172),
            .DOUT(N__6171),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__6173),
            .PADOUT(N__6172),
            .PADIN(N__6171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__6164),
            .DIN(N__6163),
            .DOUT(N__6162),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__6164),
            .PADOUT(N__6163),
            .PADIN(N__6162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5758),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_6_iopad (
            .OE(N__6155),
            .DIN(N__6154),
            .DOUT(N__6153),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__6155),
            .PADOUT(N__6154),
            .PADIN(N__6153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2740),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_serial_data_ibuf_iopad (
            .OE(N__6146),
            .DIN(N__6145),
            .DOUT(N__6144),
            .PACKAGEPIN(i_serial_data));
    defparam i_serial_data_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_serial_data_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_serial_data_ibuf_preio (
            .PADOEN(N__6146),
            .PADOUT(N__6145),
            .PADIN(N__6144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(test1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD from_ir_ibuf_iopad (
            .OE(N__6137),
            .DIN(N__6136),
            .DOUT(N__6135),
            .PACKAGEPIN(from_ir));
    defparam from_ir_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam from_ir_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO from_ir_ibuf_preio (
            .PADOEN(N__6137),
            .PADOUT(N__6136),
            .PADIN(N__6135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(test2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__6128),
            .DIN(N__6127),
            .DOUT(N__6126),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__6128),
            .PADOUT(N__6127),
            .PADIN(N__6126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5827),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__6119),
            .DIN(N__6118),
            .DOUT(N__6117),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__6119),
            .PADOUT(N__6118),
            .PADIN(N__6117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test2_obuf_iopad (
            .OE(N__6110),
            .DIN(N__6109),
            .DOUT(N__6108),
            .PACKAGEPIN(test2));
    defparam test2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test2_obuf_preio (
            .PADOEN(N__6110),
            .PADOUT(N__6109),
            .PADIN(N__6108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3816),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_5_iopad (
            .OE(N__6101),
            .DIN(N__6100),
            .DOUT(N__6099),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__6101),
            .PADOUT(N__6100),
            .PADIN(N__6099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3595),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__6092),
            .DIN(N__6091),
            .DOUT(N__6090),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__6092),
            .PADOUT(N__6091),
            .PADIN(N__6090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1357 (
            .O(N__6073),
            .I(N__6069));
    InMux I__1356 (
            .O(N__6072),
            .I(N__6066));
    LocalMux I__1355 (
            .O(N__6069),
            .I(\uut2.stateZ0Z_6 ));
    LocalMux I__1354 (
            .O(N__6066),
            .I(\uut2.stateZ0Z_6 ));
    CascadeMux I__1353 (
            .O(N__6061),
            .I(N__6058));
    InMux I__1352 (
            .O(N__6058),
            .I(N__6055));
    LocalMux I__1351 (
            .O(N__6055),
            .I(N__6052));
    Odrv4 I__1350 (
            .O(N__6052),
            .I(\uut2.tx_dataZ0Z_4 ));
    ClkMux I__1349 (
            .O(N__6049),
            .I(N__5944));
    ClkMux I__1348 (
            .O(N__6048),
            .I(N__5944));
    ClkMux I__1347 (
            .O(N__6047),
            .I(N__5944));
    ClkMux I__1346 (
            .O(N__6046),
            .I(N__5944));
    ClkMux I__1345 (
            .O(N__6045),
            .I(N__5944));
    ClkMux I__1344 (
            .O(N__6044),
            .I(N__5944));
    ClkMux I__1343 (
            .O(N__6043),
            .I(N__5944));
    ClkMux I__1342 (
            .O(N__6042),
            .I(N__5944));
    ClkMux I__1341 (
            .O(N__6041),
            .I(N__5944));
    ClkMux I__1340 (
            .O(N__6040),
            .I(N__5944));
    ClkMux I__1339 (
            .O(N__6039),
            .I(N__5944));
    ClkMux I__1338 (
            .O(N__6038),
            .I(N__5944));
    ClkMux I__1337 (
            .O(N__6037),
            .I(N__5944));
    ClkMux I__1336 (
            .O(N__6036),
            .I(N__5944));
    ClkMux I__1335 (
            .O(N__6035),
            .I(N__5944));
    ClkMux I__1334 (
            .O(N__6034),
            .I(N__5944));
    ClkMux I__1333 (
            .O(N__6033),
            .I(N__5944));
    ClkMux I__1332 (
            .O(N__6032),
            .I(N__5944));
    ClkMux I__1331 (
            .O(N__6031),
            .I(N__5944));
    ClkMux I__1330 (
            .O(N__6030),
            .I(N__5944));
    ClkMux I__1329 (
            .O(N__6029),
            .I(N__5944));
    ClkMux I__1328 (
            .O(N__6028),
            .I(N__5944));
    ClkMux I__1327 (
            .O(N__6027),
            .I(N__5944));
    ClkMux I__1326 (
            .O(N__6026),
            .I(N__5944));
    ClkMux I__1325 (
            .O(N__6025),
            .I(N__5944));
    ClkMux I__1324 (
            .O(N__6024),
            .I(N__5944));
    ClkMux I__1323 (
            .O(N__6023),
            .I(N__5944));
    ClkMux I__1322 (
            .O(N__6022),
            .I(N__5944));
    ClkMux I__1321 (
            .O(N__6021),
            .I(N__5944));
    ClkMux I__1320 (
            .O(N__6020),
            .I(N__5944));
    ClkMux I__1319 (
            .O(N__6019),
            .I(N__5944));
    ClkMux I__1318 (
            .O(N__6018),
            .I(N__5944));
    ClkMux I__1317 (
            .O(N__6017),
            .I(N__5944));
    ClkMux I__1316 (
            .O(N__6016),
            .I(N__5944));
    ClkMux I__1315 (
            .O(N__6015),
            .I(N__5944));
    GlobalMux I__1314 (
            .O(N__5944),
            .I(N__5941));
    gio2CtrlBuf I__1313 (
            .O(N__5941),
            .I(CLKOP_g));
    CEMux I__1312 (
            .O(N__5938),
            .I(N__5920));
    CEMux I__1311 (
            .O(N__5937),
            .I(N__5920));
    CEMux I__1310 (
            .O(N__5936),
            .I(N__5920));
    CEMux I__1309 (
            .O(N__5935),
            .I(N__5920));
    CEMux I__1308 (
            .O(N__5934),
            .I(N__5920));
    CEMux I__1307 (
            .O(N__5933),
            .I(N__5920));
    GlobalMux I__1306 (
            .O(N__5920),
            .I(N__5917));
    gio2CtrlBuf I__1305 (
            .O(N__5917),
            .I(N_123_g));
    InMux I__1304 (
            .O(N__5914),
            .I(N__5911));
    LocalMux I__1303 (
            .O(N__5911),
            .I(N__5897));
    SRMux I__1302 (
            .O(N__5910),
            .I(N__5854));
    SRMux I__1301 (
            .O(N__5909),
            .I(N__5854));
    SRMux I__1300 (
            .O(N__5908),
            .I(N__5854));
    SRMux I__1299 (
            .O(N__5907),
            .I(N__5854));
    SRMux I__1298 (
            .O(N__5906),
            .I(N__5854));
    SRMux I__1297 (
            .O(N__5905),
            .I(N__5854));
    SRMux I__1296 (
            .O(N__5904),
            .I(N__5854));
    SRMux I__1295 (
            .O(N__5903),
            .I(N__5854));
    SRMux I__1294 (
            .O(N__5902),
            .I(N__5854));
    SRMux I__1293 (
            .O(N__5901),
            .I(N__5854));
    SRMux I__1292 (
            .O(N__5900),
            .I(N__5854));
    Glb2LocalMux I__1291 (
            .O(N__5897),
            .I(N__5854));
    SRMux I__1290 (
            .O(N__5896),
            .I(N__5854));
    SRMux I__1289 (
            .O(N__5895),
            .I(N__5854));
    SRMux I__1288 (
            .O(N__5894),
            .I(N__5854));
    SRMux I__1287 (
            .O(N__5893),
            .I(N__5854));
    SRMux I__1286 (
            .O(N__5892),
            .I(N__5854));
    SRMux I__1285 (
            .O(N__5891),
            .I(N__5854));
    GlobalMux I__1284 (
            .O(N__5854),
            .I(N__5851));
    gio2CtrlBuf I__1283 (
            .O(N__5851),
            .I(rst_count_i_g_19));
    InMux I__1282 (
            .O(N__5848),
            .I(N__5845));
    LocalMux I__1281 (
            .O(N__5845),
            .I(N__5841));
    InMux I__1280 (
            .O(N__5844),
            .I(N__5838));
    Span4Mux_v I__1279 (
            .O(N__5841),
            .I(N__5835));
    LocalMux I__1278 (
            .O(N__5838),
            .I(N__5832));
    Odrv4 I__1277 (
            .O(N__5835),
            .I(o_rx_data_3));
    Odrv4 I__1276 (
            .O(N__5832),
            .I(o_rx_data_3));
    IoInMux I__1275 (
            .O(N__5827),
            .I(N__5824));
    LocalMux I__1274 (
            .O(N__5824),
            .I(N__5821));
    Span4Mux_s1_h I__1273 (
            .O(N__5821),
            .I(N__5818));
    Span4Mux_v I__1272 (
            .O(N__5818),
            .I(N__5815));
    Odrv4 I__1271 (
            .O(N__5815),
            .I(o_rx_data_i_3));
    InMux I__1270 (
            .O(N__5812),
            .I(N__5808));
    InMux I__1269 (
            .O(N__5811),
            .I(N__5805));
    LocalMux I__1268 (
            .O(N__5808),
            .I(N__5802));
    LocalMux I__1267 (
            .O(N__5805),
            .I(N__5799));
    Span4Mux_s2_h I__1266 (
            .O(N__5802),
            .I(N__5796));
    Odrv12 I__1265 (
            .O(N__5799),
            .I(o_rx_data_4));
    Odrv4 I__1264 (
            .O(N__5796),
            .I(o_rx_data_4));
    IoInMux I__1263 (
            .O(N__5791),
            .I(N__5788));
    LocalMux I__1262 (
            .O(N__5788),
            .I(N__5785));
    Span4Mux_s0_h I__1261 (
            .O(N__5785),
            .I(N__5782));
    Odrv4 I__1260 (
            .O(N__5782),
            .I(o_rx_data_i_4));
    InMux I__1259 (
            .O(N__5779),
            .I(N__5776));
    LocalMux I__1258 (
            .O(N__5776),
            .I(N__5772));
    InMux I__1257 (
            .O(N__5775),
            .I(N__5769));
    Span4Mux_v I__1256 (
            .O(N__5772),
            .I(N__5766));
    LocalMux I__1255 (
            .O(N__5769),
            .I(N__5763));
    Odrv4 I__1254 (
            .O(N__5766),
            .I(o_rx_data_1));
    Odrv4 I__1253 (
            .O(N__5763),
            .I(o_rx_data_1));
    IoInMux I__1252 (
            .O(N__5758),
            .I(N__5755));
    LocalMux I__1251 (
            .O(N__5755),
            .I(N__5752));
    Span4Mux_s0_h I__1250 (
            .O(N__5752),
            .I(N__5749));
    Odrv4 I__1249 (
            .O(N__5749),
            .I(o_rx_data_i_1));
    InMux I__1248 (
            .O(N__5746),
            .I(N__5743));
    LocalMux I__1247 (
            .O(N__5743),
            .I(N__5740));
    Span4Mux_v I__1246 (
            .O(N__5740),
            .I(N__5736));
    InMux I__1245 (
            .O(N__5739),
            .I(N__5733));
    Span4Mux_v I__1244 (
            .O(N__5736),
            .I(N__5730));
    LocalMux I__1243 (
            .O(N__5733),
            .I(N__5727));
    Odrv4 I__1242 (
            .O(N__5730),
            .I(o_rx_data_2));
    Odrv4 I__1241 (
            .O(N__5727),
            .I(o_rx_data_2));
    IoInMux I__1240 (
            .O(N__5722),
            .I(N__5719));
    LocalMux I__1239 (
            .O(N__5719),
            .I(o_rx_data_i_2));
    InMux I__1238 (
            .O(N__5716),
            .I(N__5712));
    InMux I__1237 (
            .O(N__5715),
            .I(N__5709));
    LocalMux I__1236 (
            .O(N__5712),
            .I(N__5706));
    LocalMux I__1235 (
            .O(N__5709),
            .I(N__5703));
    Span4Mux_v I__1234 (
            .O(N__5706),
            .I(N__5700));
    Span12Mux_s3_h I__1233 (
            .O(N__5703),
            .I(N__5697));
    Odrv4 I__1232 (
            .O(N__5700),
            .I(o_rx_data_0));
    Odrv12 I__1231 (
            .O(N__5697),
            .I(o_rx_data_0));
    IoInMux I__1230 (
            .O(N__5692),
            .I(N__5689));
    LocalMux I__1229 (
            .O(N__5689),
            .I(o_rx_data_i_0));
    InMux I__1228 (
            .O(N__5686),
            .I(N__5682));
    InMux I__1227 (
            .O(N__5685),
            .I(N__5679));
    LocalMux I__1226 (
            .O(N__5682),
            .I(\uut2.stateZ0Z_4 ));
    LocalMux I__1225 (
            .O(N__5679),
            .I(\uut2.stateZ0Z_4 ));
    CascadeMux I__1224 (
            .O(N__5674),
            .I(N__5671));
    InMux I__1223 (
            .O(N__5671),
            .I(N__5668));
    LocalMux I__1222 (
            .O(N__5668),
            .I(\uut2.serial_data_24_iv_4 ));
    InMux I__1221 (
            .O(N__5665),
            .I(N__5661));
    InMux I__1220 (
            .O(N__5664),
            .I(N__5658));
    LocalMux I__1219 (
            .O(N__5661),
            .I(N__5655));
    LocalMux I__1218 (
            .O(N__5658),
            .I(N__5652));
    Span4Mux_v I__1217 (
            .O(N__5655),
            .I(N__5649));
    Span4Mux_s2_h I__1216 (
            .O(N__5652),
            .I(N__5646));
    Odrv4 I__1215 (
            .O(N__5649),
            .I(o_rx_data_5));
    Odrv4 I__1214 (
            .O(N__5646),
            .I(o_rx_data_5));
    InMux I__1213 (
            .O(N__5641),
            .I(N__5638));
    LocalMux I__1212 (
            .O(N__5638),
            .I(\uut2.tx_dataZ0Z_5 ));
    CascadeMux I__1211 (
            .O(N__5635),
            .I(N__5632));
    InMux I__1210 (
            .O(N__5632),
            .I(N__5629));
    LocalMux I__1209 (
            .O(N__5629),
            .I(\uut2.tx_dataZ0Z_1 ));
    InMux I__1208 (
            .O(N__5626),
            .I(N__5623));
    LocalMux I__1207 (
            .O(N__5623),
            .I(\uut2.tx_dataZ0Z_0 ));
    InMux I__1206 (
            .O(N__5620),
            .I(N__5617));
    LocalMux I__1205 (
            .O(N__5617),
            .I(\uut2.tx_dataZ0Z_3 ));
    InMux I__1204 (
            .O(N__5614),
            .I(N__5611));
    LocalMux I__1203 (
            .O(N__5611),
            .I(N__5607));
    InMux I__1202 (
            .O(N__5610),
            .I(N__5604));
    Odrv4 I__1201 (
            .O(N__5607),
            .I(\uut2.stateZ0Z_8 ));
    LocalMux I__1200 (
            .O(N__5604),
            .I(\uut2.stateZ0Z_8 ));
    InMux I__1199 (
            .O(N__5599),
            .I(N__5595));
    InMux I__1198 (
            .O(N__5598),
            .I(N__5592));
    LocalMux I__1197 (
            .O(N__5595),
            .I(\uut2.stateZ0Z_7 ));
    LocalMux I__1196 (
            .O(N__5592),
            .I(\uut2.stateZ0Z_7 ));
    CascadeMux I__1195 (
            .O(N__5587),
            .I(N__5584));
    InMux I__1194 (
            .O(N__5584),
            .I(N__5581));
    LocalMux I__1193 (
            .O(N__5581),
            .I(\uut2.tx_dataZ0Z_2 ));
    InMux I__1192 (
            .O(N__5578),
            .I(N__5575));
    LocalMux I__1191 (
            .O(N__5575),
            .I(N__5571));
    InMux I__1190 (
            .O(N__5574),
            .I(N__5568));
    Odrv4 I__1189 (
            .O(N__5571),
            .I(\uut2.stateZ0Z_5 ));
    LocalMux I__1188 (
            .O(N__5568),
            .I(\uut2.stateZ0Z_5 ));
    InMux I__1187 (
            .O(N__5563),
            .I(N__5560));
    LocalMux I__1186 (
            .O(N__5560),
            .I(\uut2.serial_data_24_iv_3 ));
    InMux I__1185 (
            .O(N__5557),
            .I(N__5553));
    InMux I__1184 (
            .O(N__5556),
            .I(N__5550));
    LocalMux I__1183 (
            .O(N__5553),
            .I(N__5547));
    LocalMux I__1182 (
            .O(N__5550),
            .I(N__5544));
    Span4Mux_s3_h I__1181 (
            .O(N__5547),
            .I(N__5541));
    Odrv12 I__1180 (
            .O(N__5544),
            .I(o_rx_data_6));
    Odrv4 I__1179 (
            .O(N__5541),
            .I(o_rx_data_6));
    CascadeMux I__1178 (
            .O(N__5536),
            .I(N__5533));
    InMux I__1177 (
            .O(N__5533),
            .I(N__5530));
    LocalMux I__1176 (
            .O(N__5530),
            .I(\uut2.tx_dataZ0Z_6 ));
    InMux I__1175 (
            .O(N__5527),
            .I(N__5524));
    LocalMux I__1174 (
            .O(N__5524),
            .I(\uut2.stateZ0Z_10 ));
    InMux I__1173 (
            .O(N__5521),
            .I(N__5517));
    InMux I__1172 (
            .O(N__5520),
            .I(N__5514));
    LocalMux I__1171 (
            .O(N__5517),
            .I(\uut2.stateZ0Z_2 ));
    LocalMux I__1170 (
            .O(N__5514),
            .I(\uut2.stateZ0Z_2 ));
    InMux I__1169 (
            .O(N__5509),
            .I(N__5505));
    InMux I__1168 (
            .O(N__5508),
            .I(N__5502));
    LocalMux I__1167 (
            .O(N__5505),
            .I(\uut2.stateZ0Z_1 ));
    LocalMux I__1166 (
            .O(N__5502),
            .I(\uut2.stateZ0Z_1 ));
    InMux I__1165 (
            .O(N__5497),
            .I(N__5494));
    LocalMux I__1164 (
            .O(N__5494),
            .I(\uut2.serial_data_24_iv_2 ));
    InMux I__1163 (
            .O(N__5491),
            .I(N__5487));
    InMux I__1162 (
            .O(N__5490),
            .I(N__5484));
    LocalMux I__1161 (
            .O(N__5487),
            .I(\uut2.stateZ0Z_13 ));
    LocalMux I__1160 (
            .O(N__5484),
            .I(\uut2.stateZ0Z_13 ));
    InMux I__1159 (
            .O(N__5479),
            .I(N__5475));
    InMux I__1158 (
            .O(N__5478),
            .I(N__5472));
    LocalMux I__1157 (
            .O(N__5475),
            .I(\uut2.stateZ0Z_3 ));
    LocalMux I__1156 (
            .O(N__5472),
            .I(\uut2.stateZ0Z_3 ));
    InMux I__1155 (
            .O(N__5467),
            .I(N__5464));
    LocalMux I__1154 (
            .O(N__5464),
            .I(\uut2.serial_data_24_iv_1 ));
    InMux I__1153 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__1152 (
            .O(N__5458),
            .I(N__5455));
    Odrv12 I__1151 (
            .O(N__5455),
            .I(\uut1.rx_sampling_clockZ0 ));
    InMux I__1150 (
            .O(N__5452),
            .I(N__5448));
    InMux I__1149 (
            .O(N__5451),
            .I(N__5442));
    LocalMux I__1148 (
            .O(N__5448),
            .I(N__5439));
    InMux I__1147 (
            .O(N__5447),
            .I(N__5434));
    InMux I__1146 (
            .O(N__5446),
            .I(N__5434));
    InMux I__1145 (
            .O(N__5445),
            .I(N__5431));
    LocalMux I__1144 (
            .O(N__5442),
            .I(\uut1.rx_sampling_clock_regZ0Z1 ));
    Odrv4 I__1143 (
            .O(N__5439),
            .I(\uut1.rx_sampling_clock_regZ0Z1 ));
    LocalMux I__1142 (
            .O(N__5434),
            .I(\uut1.rx_sampling_clock_regZ0Z1 ));
    LocalMux I__1141 (
            .O(N__5431),
            .I(\uut1.rx_sampling_clock_regZ0Z1 ));
    InMux I__1140 (
            .O(N__5422),
            .I(N__5419));
    LocalMux I__1139 (
            .O(N__5419),
            .I(N__5410));
    InMux I__1138 (
            .O(N__5418),
            .I(N__5403));
    InMux I__1137 (
            .O(N__5417),
            .I(N__5403));
    InMux I__1136 (
            .O(N__5416),
            .I(N__5403));
    CascadeMux I__1135 (
            .O(N__5415),
            .I(N__5398));
    CascadeMux I__1134 (
            .O(N__5414),
            .I(N__5395));
    InMux I__1133 (
            .O(N__5413),
            .I(N__5392));
    Span4Mux_v I__1132 (
            .O(N__5410),
            .I(N__5389));
    LocalMux I__1131 (
            .O(N__5403),
            .I(N__5386));
    InMux I__1130 (
            .O(N__5402),
            .I(N__5377));
    InMux I__1129 (
            .O(N__5401),
            .I(N__5377));
    InMux I__1128 (
            .O(N__5398),
            .I(N__5377));
    InMux I__1127 (
            .O(N__5395),
            .I(N__5377));
    LocalMux I__1126 (
            .O(N__5392),
            .I(\uut1.data_validationZ0 ));
    Odrv4 I__1125 (
            .O(N__5389),
            .I(\uut1.data_validationZ0 ));
    Odrv12 I__1124 (
            .O(N__5386),
            .I(\uut1.data_validationZ0 ));
    LocalMux I__1123 (
            .O(N__5377),
            .I(\uut1.data_validationZ0 ));
    InMux I__1122 (
            .O(N__5368),
            .I(N__5363));
    CascadeMux I__1121 (
            .O(N__5367),
            .I(N__5360));
    InMux I__1120 (
            .O(N__5366),
            .I(N__5357));
    LocalMux I__1119 (
            .O(N__5363),
            .I(N__5354));
    InMux I__1118 (
            .O(N__5360),
            .I(N__5351));
    LocalMux I__1117 (
            .O(N__5357),
            .I(\uut1.rx_dataZ0Z_4 ));
    Odrv4 I__1116 (
            .O(N__5354),
            .I(\uut1.rx_dataZ0Z_4 ));
    LocalMux I__1115 (
            .O(N__5351),
            .I(\uut1.rx_dataZ0Z_4 ));
    CascadeMux I__1114 (
            .O(N__5344),
            .I(N__5336));
    CascadeMux I__1113 (
            .O(N__5343),
            .I(N__5333));
    InMux I__1112 (
            .O(N__5342),
            .I(N__5330));
    InMux I__1111 (
            .O(N__5341),
            .I(N__5327));
    InMux I__1110 (
            .O(N__5340),
            .I(N__5319));
    InMux I__1109 (
            .O(N__5339),
            .I(N__5319));
    InMux I__1108 (
            .O(N__5336),
            .I(N__5315));
    InMux I__1107 (
            .O(N__5333),
            .I(N__5312));
    LocalMux I__1106 (
            .O(N__5330),
            .I(N__5307));
    LocalMux I__1105 (
            .O(N__5327),
            .I(N__5307));
    InMux I__1104 (
            .O(N__5326),
            .I(N__5300));
    InMux I__1103 (
            .O(N__5325),
            .I(N__5300));
    InMux I__1102 (
            .O(N__5324),
            .I(N__5300));
    LocalMux I__1101 (
            .O(N__5319),
            .I(N__5297));
    InMux I__1100 (
            .O(N__5318),
            .I(N__5294));
    LocalMux I__1099 (
            .O(N__5315),
            .I(N__5287));
    LocalMux I__1098 (
            .O(N__5312),
            .I(N__5287));
    Span4Mux_v I__1097 (
            .O(N__5307),
            .I(N__5287));
    LocalMux I__1096 (
            .O(N__5300),
            .I(N__5284));
    Span4Mux_h I__1095 (
            .O(N__5297),
            .I(N__5279));
    LocalMux I__1094 (
            .O(N__5294),
            .I(N__5279));
    Odrv4 I__1093 (
            .O(N__5287),
            .I(\uut1.modem_serial_dataZ0 ));
    Odrv12 I__1092 (
            .O(N__5284),
            .I(\uut1.modem_serial_dataZ0 ));
    Odrv4 I__1091 (
            .O(N__5279),
            .I(\uut1.modem_serial_dataZ0 ));
    CEMux I__1090 (
            .O(N__5272),
            .I(N__5269));
    LocalMux I__1089 (
            .O(N__5269),
            .I(N__5263));
    InMux I__1088 (
            .O(N__5268),
            .I(N__5256));
    InMux I__1087 (
            .O(N__5267),
            .I(N__5256));
    InMux I__1086 (
            .O(N__5266),
            .I(N__5253));
    Span4Mux_h I__1085 (
            .O(N__5263),
            .I(N__5247));
    InMux I__1084 (
            .O(N__5262),
            .I(N__5242));
    InMux I__1083 (
            .O(N__5261),
            .I(N__5242));
    LocalMux I__1082 (
            .O(N__5256),
            .I(N__5239));
    LocalMux I__1081 (
            .O(N__5253),
            .I(N__5236));
    InMux I__1080 (
            .O(N__5252),
            .I(N__5229));
    InMux I__1079 (
            .O(N__5251),
            .I(N__5229));
    InMux I__1078 (
            .O(N__5250),
            .I(N__5229));
    Odrv4 I__1077 (
            .O(N__5247),
            .I(\uut1.rx_sample_en ));
    LocalMux I__1076 (
            .O(N__5242),
            .I(\uut1.rx_sample_en ));
    Odrv4 I__1075 (
            .O(N__5239),
            .I(\uut1.rx_sample_en ));
    Odrv4 I__1074 (
            .O(N__5236),
            .I(\uut1.rx_sample_en ));
    LocalMux I__1073 (
            .O(N__5229),
            .I(\uut1.rx_sample_en ));
    CascadeMux I__1072 (
            .O(N__5218),
            .I(N__5214));
    CascadeMux I__1071 (
            .O(N__5217),
            .I(N__5211));
    InMux I__1070 (
            .O(N__5214),
            .I(N__5207));
    InMux I__1069 (
            .O(N__5211),
            .I(N__5204));
    InMux I__1068 (
            .O(N__5210),
            .I(N__5201));
    LocalMux I__1067 (
            .O(N__5207),
            .I(N__5198));
    LocalMux I__1066 (
            .O(N__5204),
            .I(\uut1.rx_dataZ0Z_9 ));
    LocalMux I__1065 (
            .O(N__5201),
            .I(\uut1.rx_dataZ0Z_9 ));
    Odrv4 I__1064 (
            .O(N__5198),
            .I(\uut1.rx_dataZ0Z_9 ));
    InMux I__1063 (
            .O(N__5191),
            .I(N__5184));
    InMux I__1062 (
            .O(N__5190),
            .I(N__5181));
    InMux I__1061 (
            .O(N__5189),
            .I(N__5176));
    InMux I__1060 (
            .O(N__5188),
            .I(N__5173));
    InMux I__1059 (
            .O(N__5187),
            .I(N__5170));
    LocalMux I__1058 (
            .O(N__5184),
            .I(N__5165));
    LocalMux I__1057 (
            .O(N__5181),
            .I(N__5165));
    InMux I__1056 (
            .O(N__5180),
            .I(N__5162));
    InMux I__1055 (
            .O(N__5179),
            .I(N__5159));
    LocalMux I__1054 (
            .O(N__5176),
            .I(\uut1.stateZ0Z_2 ));
    LocalMux I__1053 (
            .O(N__5173),
            .I(\uut1.stateZ0Z_2 ));
    LocalMux I__1052 (
            .O(N__5170),
            .I(\uut1.stateZ0Z_2 ));
    Odrv4 I__1051 (
            .O(N__5165),
            .I(\uut1.stateZ0Z_2 ));
    LocalMux I__1050 (
            .O(N__5162),
            .I(\uut1.stateZ0Z_2 ));
    LocalMux I__1049 (
            .O(N__5159),
            .I(\uut1.stateZ0Z_2 ));
    InMux I__1048 (
            .O(N__5146),
            .I(N__5143));
    LocalMux I__1047 (
            .O(N__5143),
            .I(\uut1.rx_data_7_m_9 ));
    InMux I__1046 (
            .O(N__5140),
            .I(N__5136));
    InMux I__1045 (
            .O(N__5139),
            .I(N__5133));
    LocalMux I__1044 (
            .O(N__5136),
            .I(\uut2.stateZ0Z_11 ));
    LocalMux I__1043 (
            .O(N__5133),
            .I(\uut2.stateZ0Z_11 ));
    IoInMux I__1042 (
            .O(N__5128),
            .I(N__5124));
    CascadeMux I__1041 (
            .O(N__5127),
            .I(N__5121));
    LocalMux I__1040 (
            .O(N__5124),
            .I(N__5118));
    InMux I__1039 (
            .O(N__5121),
            .I(N__5115));
    Span12Mux_s4_h I__1038 (
            .O(N__5118),
            .I(N__5112));
    LocalMux I__1037 (
            .O(N__5115),
            .I(N__5109));
    Odrv12 I__1036 (
            .O(N__5112),
            .I(count_RNIH42R1Z0Z_2));
    Odrv4 I__1035 (
            .O(N__5109),
            .I(count_RNIH42R1Z0Z_2));
    InMux I__1034 (
            .O(N__5104),
            .I(N__5095));
    InMux I__1033 (
            .O(N__5103),
            .I(N__5095));
    InMux I__1032 (
            .O(N__5102),
            .I(N__5095));
    LocalMux I__1031 (
            .O(N__5095),
            .I(N__5092));
    Span4Mux_s3_h I__1030 (
            .O(N__5092),
            .I(N__5089));
    Odrv4 I__1029 (
            .O(N__5089),
            .I(i_start_tx_0));
    CascadeMux I__1028 (
            .O(N__5086),
            .I(N__5083));
    InMux I__1027 (
            .O(N__5083),
            .I(N__5074));
    InMux I__1026 (
            .O(N__5082),
            .I(N__5074));
    InMux I__1025 (
            .O(N__5081),
            .I(N__5074));
    LocalMux I__1024 (
            .O(N__5074),
            .I(\uut2.stateZ0Z_0 ));
    IoInMux I__1023 (
            .O(N__5071),
            .I(N__5068));
    LocalMux I__1022 (
            .O(N__5068),
            .I(N__5065));
    Span12Mux_s10_h I__1021 (
            .O(N__5065),
            .I(N__5062));
    Odrv12 I__1020 (
            .O(N__5062),
            .I(o_serial_data_c));
    CEMux I__1019 (
            .O(N__5059),
            .I(N__5056));
    LocalMux I__1018 (
            .O(N__5056),
            .I(N__5053));
    Span4Mux_s1_h I__1017 (
            .O(N__5053),
            .I(N__5050));
    Odrv4 I__1016 (
            .O(N__5050),
            .I(\uut2.serial_data_RNOZ0Z_0 ));
    InMux I__1015 (
            .O(N__5047),
            .I(N__5042));
    InMux I__1014 (
            .O(N__5046),
            .I(N__5038));
    InMux I__1013 (
            .O(N__5045),
            .I(N__5035));
    LocalMux I__1012 (
            .O(N__5042),
            .I(N__5032));
    InMux I__1011 (
            .O(N__5041),
            .I(N__5029));
    LocalMux I__1010 (
            .O(N__5038),
            .I(\uut1.stateZ0Z_1 ));
    LocalMux I__1009 (
            .O(N__5035),
            .I(\uut1.stateZ0Z_1 ));
    Odrv4 I__1008 (
            .O(N__5032),
            .I(\uut1.stateZ0Z_1 ));
    LocalMux I__1007 (
            .O(N__5029),
            .I(\uut1.stateZ0Z_1 ));
    InMux I__1006 (
            .O(N__5020),
            .I(N__5011));
    InMux I__1005 (
            .O(N__5019),
            .I(N__5011));
    CascadeMux I__1004 (
            .O(N__5018),
            .I(N__5008));
    CascadeMux I__1003 (
            .O(N__5017),
            .I(N__5004));
    InMux I__1002 (
            .O(N__5016),
            .I(N__5000));
    LocalMux I__1001 (
            .O(N__5011),
            .I(N__4997));
    InMux I__1000 (
            .O(N__5008),
            .I(N__4994));
    InMux I__999 (
            .O(N__5007),
            .I(N__4991));
    InMux I__998 (
            .O(N__5004),
            .I(N__4988));
    InMux I__997 (
            .O(N__5003),
            .I(N__4985));
    LocalMux I__996 (
            .O(N__5000),
            .I(\uut1.stateZ0Z_11 ));
    Odrv4 I__995 (
            .O(N__4997),
            .I(\uut1.stateZ0Z_11 ));
    LocalMux I__994 (
            .O(N__4994),
            .I(\uut1.stateZ0Z_11 ));
    LocalMux I__993 (
            .O(N__4991),
            .I(\uut1.stateZ0Z_11 ));
    LocalMux I__992 (
            .O(N__4988),
            .I(\uut1.stateZ0Z_11 ));
    LocalMux I__991 (
            .O(N__4985),
            .I(\uut1.stateZ0Z_11 ));
    InMux I__990 (
            .O(N__4972),
            .I(N__4966));
    InMux I__989 (
            .O(N__4971),
            .I(N__4963));
    InMux I__988 (
            .O(N__4970),
            .I(N__4959));
    InMux I__987 (
            .O(N__4969),
            .I(N__4956));
    LocalMux I__986 (
            .O(N__4966),
            .I(N__4951));
    LocalMux I__985 (
            .O(N__4963),
            .I(N__4951));
    InMux I__984 (
            .O(N__4962),
            .I(N__4948));
    LocalMux I__983 (
            .O(N__4959),
            .I(\uut1.stateZ0Z_0 ));
    LocalMux I__982 (
            .O(N__4956),
            .I(\uut1.stateZ0Z_0 ));
    Odrv4 I__981 (
            .O(N__4951),
            .I(\uut1.stateZ0Z_0 ));
    LocalMux I__980 (
            .O(N__4948),
            .I(\uut1.stateZ0Z_0 ));
    CascadeMux I__979 (
            .O(N__4939),
            .I(\uut1.rx_sample_en_cascade_ ));
    InMux I__978 (
            .O(N__4936),
            .I(N__4932));
    InMux I__977 (
            .O(N__4935),
            .I(N__4925));
    LocalMux I__976 (
            .O(N__4932),
            .I(N__4922));
    InMux I__975 (
            .O(N__4931),
            .I(N__4919));
    InMux I__974 (
            .O(N__4930),
            .I(N__4916));
    InMux I__973 (
            .O(N__4929),
            .I(N__4913));
    InMux I__972 (
            .O(N__4928),
            .I(N__4910));
    LocalMux I__971 (
            .O(N__4925),
            .I(\uut1.stateZ0Z_3 ));
    Odrv4 I__970 (
            .O(N__4922),
            .I(\uut1.stateZ0Z_3 ));
    LocalMux I__969 (
            .O(N__4919),
            .I(\uut1.stateZ0Z_3 ));
    LocalMux I__968 (
            .O(N__4916),
            .I(\uut1.stateZ0Z_3 ));
    LocalMux I__967 (
            .O(N__4913),
            .I(\uut1.stateZ0Z_3 ));
    LocalMux I__966 (
            .O(N__4910),
            .I(\uut1.stateZ0Z_3 ));
    CascadeMux I__965 (
            .O(N__4897),
            .I(\uut1.rx_data_10_m_8_cascade_ ));
    InMux I__964 (
            .O(N__4894),
            .I(N__4891));
    LocalMux I__963 (
            .O(N__4891),
            .I(\uut1.N_220_0 ));
    InMux I__962 (
            .O(N__4888),
            .I(N__4883));
    InMux I__961 (
            .O(N__4887),
            .I(N__4878));
    InMux I__960 (
            .O(N__4886),
            .I(N__4878));
    LocalMux I__959 (
            .O(N__4883),
            .I(\uut1.rx_dataZ0Z_8 ));
    LocalMux I__958 (
            .O(N__4878),
            .I(\uut1.rx_dataZ0Z_8 ));
    InMux I__957 (
            .O(N__4873),
            .I(N__4869));
    CascadeMux I__956 (
            .O(N__4872),
            .I(N__4865));
    LocalMux I__955 (
            .O(N__4869),
            .I(N__4861));
    InMux I__954 (
            .O(N__4868),
            .I(N__4856));
    InMux I__953 (
            .O(N__4865),
            .I(N__4856));
    InMux I__952 (
            .O(N__4864),
            .I(N__4853));
    Odrv4 I__951 (
            .O(N__4861),
            .I(\uut1.rx_sampling_clock_regZ0Z2 ));
    LocalMux I__950 (
            .O(N__4856),
            .I(\uut1.rx_sampling_clock_regZ0Z2 ));
    LocalMux I__949 (
            .O(N__4853),
            .I(\uut1.rx_sampling_clock_regZ0Z2 ));
    InMux I__948 (
            .O(N__4846),
            .I(N__4837));
    InMux I__947 (
            .O(N__4845),
            .I(N__4832));
    InMux I__946 (
            .O(N__4844),
            .I(N__4832));
    InMux I__945 (
            .O(N__4843),
            .I(N__4829));
    InMux I__944 (
            .O(N__4842),
            .I(N__4826));
    InMux I__943 (
            .O(N__4841),
            .I(N__4821));
    InMux I__942 (
            .O(N__4840),
            .I(N__4821));
    LocalMux I__941 (
            .O(N__4837),
            .I(\uut1.state_RNID38FZ0Z_1 ));
    LocalMux I__940 (
            .O(N__4832),
            .I(\uut1.state_RNID38FZ0Z_1 ));
    LocalMux I__939 (
            .O(N__4829),
            .I(\uut1.state_RNID38FZ0Z_1 ));
    LocalMux I__938 (
            .O(N__4826),
            .I(\uut1.state_RNID38FZ0Z_1 ));
    LocalMux I__937 (
            .O(N__4821),
            .I(\uut1.state_RNID38FZ0Z_1 ));
    InMux I__936 (
            .O(N__4810),
            .I(N__4807));
    LocalMux I__935 (
            .O(N__4807),
            .I(\uut1.N_221_0 ));
    CascadeMux I__934 (
            .O(N__4804),
            .I(N__4800));
    CascadeMux I__933 (
            .O(N__4803),
            .I(N__4797));
    InMux I__932 (
            .O(N__4800),
            .I(N__4793));
    InMux I__931 (
            .O(N__4797),
            .I(N__4790));
    InMux I__930 (
            .O(N__4796),
            .I(N__4787));
    LocalMux I__929 (
            .O(N__4793),
            .I(N__4784));
    LocalMux I__928 (
            .O(N__4790),
            .I(\uut1.rx_dataZ0Z_5 ));
    LocalMux I__927 (
            .O(N__4787),
            .I(\uut1.rx_dataZ0Z_5 ));
    Odrv4 I__926 (
            .O(N__4784),
            .I(\uut1.rx_dataZ0Z_5 ));
    CascadeMux I__925 (
            .O(N__4777),
            .I(\uut1.rx_sampling_counter16_cascade_ ));
    InMux I__924 (
            .O(N__4774),
            .I(N__4766));
    InMux I__923 (
            .O(N__4773),
            .I(N__4766));
    InMux I__922 (
            .O(N__4772),
            .I(N__4761));
    InMux I__921 (
            .O(N__4771),
            .I(N__4761));
    LocalMux I__920 (
            .O(N__4766),
            .I(\uut1.rx_sampling_counter_1_sqmuxa ));
    LocalMux I__919 (
            .O(N__4761),
            .I(\uut1.rx_sampling_counter_1_sqmuxa ));
    InMux I__918 (
            .O(N__4756),
            .I(N__4750));
    InMux I__917 (
            .O(N__4755),
            .I(N__4747));
    InMux I__916 (
            .O(N__4754),
            .I(N__4742));
    InMux I__915 (
            .O(N__4753),
            .I(N__4742));
    LocalMux I__914 (
            .O(N__4750),
            .I(clk_countZ0Z_0));
    LocalMux I__913 (
            .O(N__4747),
            .I(clk_countZ0Z_0));
    LocalMux I__912 (
            .O(N__4742),
            .I(clk_countZ0Z_0));
    InMux I__911 (
            .O(N__4735),
            .I(N__4730));
    InMux I__910 (
            .O(N__4734),
            .I(N__4727));
    InMux I__909 (
            .O(N__4733),
            .I(N__4724));
    LocalMux I__908 (
            .O(N__4730),
            .I(\uut1.rx_sampling_startZ0 ));
    LocalMux I__907 (
            .O(N__4727),
            .I(\uut1.rx_sampling_startZ0 ));
    LocalMux I__906 (
            .O(N__4724),
            .I(\uut1.rx_sampling_startZ0 ));
    InMux I__905 (
            .O(N__4717),
            .I(N__4713));
    InMux I__904 (
            .O(N__4716),
            .I(N__4710));
    LocalMux I__903 (
            .O(N__4713),
            .I(N__4707));
    LocalMux I__902 (
            .O(N__4710),
            .I(N__4702));
    Span4Mux_h I__901 (
            .O(N__4707),
            .I(N__4702));
    Odrv4 I__900 (
            .O(N__4702),
            .I(\uut1.rx_data_ready_regZ0Z1 ));
    InMux I__899 (
            .O(N__4699),
            .I(N__4696));
    LocalMux I__898 (
            .O(N__4696),
            .I(N__4693));
    Span4Mux_h I__897 (
            .O(N__4693),
            .I(N__4690));
    Odrv4 I__896 (
            .O(N__4690),
            .I(\uut1.rx_data_ready_regZ0Z2 ));
    CascadeMux I__895 (
            .O(N__4687),
            .I(N__4682));
    InMux I__894 (
            .O(N__4686),
            .I(N__4679));
    CascadeMux I__893 (
            .O(N__4685),
            .I(N__4676));
    InMux I__892 (
            .O(N__4682),
            .I(N__4673));
    LocalMux I__891 (
            .O(N__4679),
            .I(N__4670));
    InMux I__890 (
            .O(N__4676),
            .I(N__4667));
    LocalMux I__889 (
            .O(N__4673),
            .I(\uut1.rx_dataZ0Z_7 ));
    Odrv4 I__888 (
            .O(N__4670),
            .I(\uut1.rx_dataZ0Z_7 ));
    LocalMux I__887 (
            .O(N__4667),
            .I(\uut1.rx_dataZ0Z_7 ));
    CascadeMux I__886 (
            .O(N__4660),
            .I(N__4657));
    InMux I__885 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__884 (
            .O(N__4654),
            .I(N__4650));
    InMux I__883 (
            .O(N__4653),
            .I(N__4647));
    Odrv4 I__882 (
            .O(N__4650),
            .I(\uut1.state_ns_a2_0_0_2 ));
    LocalMux I__881 (
            .O(N__4647),
            .I(\uut1.state_ns_a2_0_0_2 ));
    InMux I__880 (
            .O(N__4642),
            .I(N__4637));
    InMux I__879 (
            .O(N__4641),
            .I(N__4634));
    CascadeMux I__878 (
            .O(N__4640),
            .I(N__4631));
    LocalMux I__877 (
            .O(N__4637),
            .I(N__4626));
    LocalMux I__876 (
            .O(N__4634),
            .I(N__4626));
    InMux I__875 (
            .O(N__4631),
            .I(N__4623));
    Odrv12 I__874 (
            .O(N__4626),
            .I(\uut1.rx_dataZ0Z_6 ));
    LocalMux I__873 (
            .O(N__4623),
            .I(\uut1.rx_dataZ0Z_6 ));
    InMux I__872 (
            .O(N__4618),
            .I(N__4615));
    LocalMux I__871 (
            .O(N__4615),
            .I(\uut1.rx_data_25_m_3 ));
    InMux I__870 (
            .O(N__4612),
            .I(N__4609));
    LocalMux I__869 (
            .O(N__4609),
            .I(\uut1.N_215_0 ));
    InMux I__868 (
            .O(N__4606),
            .I(N__4603));
    LocalMux I__867 (
            .O(N__4603),
            .I(\uut1.rx_data_19_m_5 ));
    CascadeMux I__866 (
            .O(N__4600),
            .I(N__4596));
    CascadeMux I__865 (
            .O(N__4599),
            .I(N__4593));
    InMux I__864 (
            .O(N__4596),
            .I(N__4589));
    InMux I__863 (
            .O(N__4593),
            .I(N__4584));
    InMux I__862 (
            .O(N__4592),
            .I(N__4584));
    LocalMux I__861 (
            .O(N__4589),
            .I(N__4581));
    LocalMux I__860 (
            .O(N__4584),
            .I(\uut1.rx_dataZ0Z_3 ));
    Odrv4 I__859 (
            .O(N__4581),
            .I(\uut1.rx_dataZ0Z_3 ));
    InMux I__858 (
            .O(N__4576),
            .I(N__4571));
    InMux I__857 (
            .O(N__4575),
            .I(N__4566));
    InMux I__856 (
            .O(N__4574),
            .I(N__4563));
    LocalMux I__855 (
            .O(N__4571),
            .I(N__4560));
    InMux I__854 (
            .O(N__4570),
            .I(N__4555));
    InMux I__853 (
            .O(N__4569),
            .I(N__4555));
    LocalMux I__852 (
            .O(N__4566),
            .I(\uut1.stateZ0Z_8 ));
    LocalMux I__851 (
            .O(N__4563),
            .I(\uut1.stateZ0Z_8 ));
    Odrv4 I__850 (
            .O(N__4560),
            .I(\uut1.stateZ0Z_8 ));
    LocalMux I__849 (
            .O(N__4555),
            .I(\uut1.stateZ0Z_8 ));
    InMux I__848 (
            .O(N__4546),
            .I(N__4542));
    InMux I__847 (
            .O(N__4545),
            .I(N__4536));
    LocalMux I__846 (
            .O(N__4542),
            .I(N__4533));
    InMux I__845 (
            .O(N__4541),
            .I(N__4530));
    InMux I__844 (
            .O(N__4540),
            .I(N__4525));
    InMux I__843 (
            .O(N__4539),
            .I(N__4525));
    LocalMux I__842 (
            .O(N__4536),
            .I(\uut1.stateZ0Z_7 ));
    Odrv4 I__841 (
            .O(N__4533),
            .I(\uut1.stateZ0Z_7 ));
    LocalMux I__840 (
            .O(N__4530),
            .I(\uut1.stateZ0Z_7 ));
    LocalMux I__839 (
            .O(N__4525),
            .I(\uut1.stateZ0Z_7 ));
    InMux I__838 (
            .O(N__4516),
            .I(N__4512));
    InMux I__837 (
            .O(N__4515),
            .I(N__4509));
    LocalMux I__836 (
            .O(N__4512),
            .I(\uut1.N_217_0_4 ));
    LocalMux I__835 (
            .O(N__4509),
            .I(\uut1.N_217_0_4 ));
    InMux I__834 (
            .O(N__4504),
            .I(N__4501));
    LocalMux I__833 (
            .O(N__4501),
            .I(\uut1.N_217_0 ));
    CEMux I__832 (
            .O(N__4498),
            .I(N__4495));
    LocalMux I__831 (
            .O(N__4495),
            .I(N__4492));
    Span4Mux_s2_v I__830 (
            .O(N__4492),
            .I(N__4489));
    Span4Mux_s2_h I__829 (
            .O(N__4489),
            .I(N__4486));
    Odrv4 I__828 (
            .O(N__4486),
            .I(\uut1.rx_sampling_clock_RNOZ0 ));
    CascadeMux I__827 (
            .O(N__4483),
            .I(N__4480));
    InMux I__826 (
            .O(N__4480),
            .I(N__4477));
    LocalMux I__825 (
            .O(N__4477),
            .I(\uut1.CO2 ));
    CascadeMux I__824 (
            .O(N__4474),
            .I(N__4471));
    InMux I__823 (
            .O(N__4471),
            .I(N__4468));
    LocalMux I__822 (
            .O(N__4468),
            .I(\uut1.N_5 ));
    InMux I__821 (
            .O(N__4465),
            .I(N__4459));
    InMux I__820 (
            .O(N__4464),
            .I(N__4452));
    InMux I__819 (
            .O(N__4463),
            .I(N__4452));
    InMux I__818 (
            .O(N__4462),
            .I(N__4452));
    LocalMux I__817 (
            .O(N__4459),
            .I(\uut1.rx_sampling_counterZ0Z_2 ));
    LocalMux I__816 (
            .O(N__4452),
            .I(\uut1.rx_sampling_counterZ0Z_2 ));
    CascadeMux I__815 (
            .O(N__4447),
            .I(N__4444));
    InMux I__814 (
            .O(N__4444),
            .I(N__4438));
    InMux I__813 (
            .O(N__4443),
            .I(N__4433));
    InMux I__812 (
            .O(N__4442),
            .I(N__4433));
    InMux I__811 (
            .O(N__4441),
            .I(N__4430));
    LocalMux I__810 (
            .O(N__4438),
            .I(\uut1.rx_sampling_counterZ0Z_1 ));
    LocalMux I__809 (
            .O(N__4433),
            .I(\uut1.rx_sampling_counterZ0Z_1 ));
    LocalMux I__808 (
            .O(N__4430),
            .I(\uut1.rx_sampling_counterZ0Z_1 ));
    CascadeMux I__807 (
            .O(N__4423),
            .I(N__4418));
    InMux I__806 (
            .O(N__4422),
            .I(N__4415));
    InMux I__805 (
            .O(N__4421),
            .I(N__4412));
    InMux I__804 (
            .O(N__4418),
            .I(N__4409));
    LocalMux I__803 (
            .O(N__4415),
            .I(\uut1.rx_sampling_counterZ0Z_3 ));
    LocalMux I__802 (
            .O(N__4412),
            .I(\uut1.rx_sampling_counterZ0Z_3 ));
    LocalMux I__801 (
            .O(N__4409),
            .I(\uut1.rx_sampling_counterZ0Z_3 ));
    InMux I__800 (
            .O(N__4402),
            .I(N__4393));
    InMux I__799 (
            .O(N__4401),
            .I(N__4393));
    InMux I__798 (
            .O(N__4400),
            .I(N__4386));
    InMux I__797 (
            .O(N__4399),
            .I(N__4386));
    InMux I__796 (
            .O(N__4398),
            .I(N__4386));
    LocalMux I__795 (
            .O(N__4393),
            .I(\uut1.rx_sampling_counterZ0Z_0 ));
    LocalMux I__794 (
            .O(N__4386),
            .I(\uut1.rx_sampling_counterZ0Z_0 ));
    InMux I__793 (
            .O(N__4381),
            .I(N__4378));
    LocalMux I__792 (
            .O(N__4378),
            .I(\uut1.rx_data_22_m_4 ));
    CascadeMux I__791 (
            .O(N__4375),
            .I(\uut1.N_221_0_5_cascade_ ));
    InMux I__790 (
            .O(N__4372),
            .I(N__4367));
    InMux I__789 (
            .O(N__4371),
            .I(N__4364));
    InMux I__788 (
            .O(N__4370),
            .I(N__4361));
    LocalMux I__787 (
            .O(N__4367),
            .I(\uut1.N_221_0_5 ));
    LocalMux I__786 (
            .O(N__4364),
            .I(\uut1.N_221_0_5 ));
    LocalMux I__785 (
            .O(N__4361),
            .I(\uut1.N_221_0_5 ));
    CascadeMux I__784 (
            .O(N__4354),
            .I(N__4348));
    CascadeMux I__783 (
            .O(N__4353),
            .I(N__4343));
    InMux I__782 (
            .O(N__4352),
            .I(N__4340));
    InMux I__781 (
            .O(N__4351),
            .I(N__4337));
    InMux I__780 (
            .O(N__4348),
            .I(N__4332));
    InMux I__779 (
            .O(N__4347),
            .I(N__4332));
    InMux I__778 (
            .O(N__4346),
            .I(N__4329));
    InMux I__777 (
            .O(N__4343),
            .I(N__4326));
    LocalMux I__776 (
            .O(N__4340),
            .I(\uut1.stateZ0Z_4 ));
    LocalMux I__775 (
            .O(N__4337),
            .I(\uut1.stateZ0Z_4 ));
    LocalMux I__774 (
            .O(N__4332),
            .I(\uut1.stateZ0Z_4 ));
    LocalMux I__773 (
            .O(N__4329),
            .I(\uut1.stateZ0Z_4 ));
    LocalMux I__772 (
            .O(N__4326),
            .I(\uut1.stateZ0Z_4 ));
    InMux I__771 (
            .O(N__4315),
            .I(N__4309));
    InMux I__770 (
            .O(N__4314),
            .I(N__4309));
    LocalMux I__769 (
            .O(N__4309),
            .I(\uut1.N_221_0_2 ));
    InMux I__768 (
            .O(N__4306),
            .I(N__4298));
    InMux I__767 (
            .O(N__4305),
            .I(N__4295));
    InMux I__766 (
            .O(N__4304),
            .I(N__4290));
    InMux I__765 (
            .O(N__4303),
            .I(N__4290));
    InMux I__764 (
            .O(N__4302),
            .I(N__4287));
    InMux I__763 (
            .O(N__4301),
            .I(N__4284));
    LocalMux I__762 (
            .O(N__4298),
            .I(\uut1.stateZ0Z_6 ));
    LocalMux I__761 (
            .O(N__4295),
            .I(\uut1.stateZ0Z_6 ));
    LocalMux I__760 (
            .O(N__4290),
            .I(\uut1.stateZ0Z_6 ));
    LocalMux I__759 (
            .O(N__4287),
            .I(\uut1.stateZ0Z_6 ));
    LocalMux I__758 (
            .O(N__4284),
            .I(\uut1.stateZ0Z_6 ));
    InMux I__757 (
            .O(N__4273),
            .I(un3_clk_count_cry_1));
    InMux I__756 (
            .O(N__4270),
            .I(un3_clk_count_cry_2));
    InMux I__755 (
            .O(N__4267),
            .I(un3_clk_count_cry_3));
    InMux I__754 (
            .O(N__4264),
            .I(un3_clk_count_cry_4));
    InMux I__753 (
            .O(N__4261),
            .I(N__4257));
    InMux I__752 (
            .O(N__4260),
            .I(N__4254));
    LocalMux I__751 (
            .O(N__4257),
            .I(clk_countZ0Z_5));
    LocalMux I__750 (
            .O(N__4254),
            .I(clk_countZ0Z_5));
    InMux I__749 (
            .O(N__4249),
            .I(N__4239));
    InMux I__748 (
            .O(N__4248),
            .I(N__4239));
    CascadeMux I__747 (
            .O(N__4247),
            .I(N__4235));
    CascadeMux I__746 (
            .O(N__4246),
            .I(N__4232));
    InMux I__745 (
            .O(N__4245),
            .I(N__4227));
    InMux I__744 (
            .O(N__4244),
            .I(N__4227));
    LocalMux I__743 (
            .O(N__4239),
            .I(N__4224));
    InMux I__742 (
            .O(N__4238),
            .I(N__4217));
    InMux I__741 (
            .O(N__4235),
            .I(N__4217));
    InMux I__740 (
            .O(N__4232),
            .I(N__4217));
    LocalMux I__739 (
            .O(N__4227),
            .I(clk_countZ0Z_2));
    Odrv4 I__738 (
            .O(N__4224),
            .I(clk_countZ0Z_2));
    LocalMux I__737 (
            .O(N__4217),
            .I(clk_countZ0Z_2));
    InMux I__736 (
            .O(N__4210),
            .I(N__4207));
    LocalMux I__735 (
            .O(N__4207),
            .I(clk_count_RNO_0Z0Z_3));
    CascadeMux I__734 (
            .O(N__4204),
            .I(N__4199));
    CascadeMux I__733 (
            .O(N__4203),
            .I(N__4196));
    InMux I__732 (
            .O(N__4202),
            .I(N__4190));
    InMux I__731 (
            .O(N__4199),
            .I(N__4190));
    InMux I__730 (
            .O(N__4196),
            .I(N__4182));
    InMux I__729 (
            .O(N__4195),
            .I(N__4182));
    LocalMux I__728 (
            .O(N__4190),
            .I(N__4179));
    InMux I__727 (
            .O(N__4189),
            .I(N__4172));
    InMux I__726 (
            .O(N__4188),
            .I(N__4172));
    InMux I__725 (
            .O(N__4187),
            .I(N__4172));
    LocalMux I__724 (
            .O(N__4182),
            .I(clk_countZ0Z_4));
    Odrv4 I__723 (
            .O(N__4179),
            .I(clk_countZ0Z_4));
    LocalMux I__722 (
            .O(N__4172),
            .I(clk_countZ0Z_4));
    InMux I__721 (
            .O(N__4165),
            .I(N__4158));
    InMux I__720 (
            .O(N__4164),
            .I(N__4153));
    InMux I__719 (
            .O(N__4163),
            .I(N__4153));
    InMux I__718 (
            .O(N__4162),
            .I(N__4148));
    InMux I__717 (
            .O(N__4161),
            .I(N__4148));
    LocalMux I__716 (
            .O(N__4158),
            .I(CLKOS3_3));
    LocalMux I__715 (
            .O(N__4153),
            .I(CLKOS3_3));
    LocalMux I__714 (
            .O(N__4148),
            .I(CLKOS3_3));
    CascadeMux I__713 (
            .O(N__4141),
            .I(N__4137));
    InMux I__712 (
            .O(N__4140),
            .I(N__4134));
    InMux I__711 (
            .O(N__4137),
            .I(N__4131));
    LocalMux I__710 (
            .O(N__4134),
            .I(clk_countZ0Z_3));
    LocalMux I__709 (
            .O(N__4131),
            .I(clk_countZ0Z_3));
    InMux I__708 (
            .O(N__4126),
            .I(N__4123));
    LocalMux I__707 (
            .O(N__4123),
            .I(\uut1.rx_data_16_m_6 ));
    InMux I__706 (
            .O(N__4120),
            .I(N__4117));
    LocalMux I__705 (
            .O(N__4117),
            .I(\uut1.rx_data_13_m_7 ));
    InMux I__704 (
            .O(N__4114),
            .I(N__4108));
    InMux I__703 (
            .O(N__4113),
            .I(N__4105));
    InMux I__702 (
            .O(N__4112),
            .I(N__4100));
    InMux I__701 (
            .O(N__4111),
            .I(N__4100));
    LocalMux I__700 (
            .O(N__4108),
            .I(\uut1.stateZ0Z_5 ));
    LocalMux I__699 (
            .O(N__4105),
            .I(\uut1.stateZ0Z_5 ));
    LocalMux I__698 (
            .O(N__4100),
            .I(\uut1.stateZ0Z_5 ));
    CascadeMux I__697 (
            .O(N__4093),
            .I(\uut1.N_221_0_2_cascade_ ));
    InMux I__696 (
            .O(N__4090),
            .I(N__4087));
    LocalMux I__695 (
            .O(N__4087),
            .I(\uut1.N_219_0 ));
    CascadeMux I__694 (
            .O(N__4084),
            .I(\uut1.rx_sampling_clock_cnv_1_cascade_ ));
    CascadeMux I__693 (
            .O(N__4081),
            .I(clk_count_RNO_0Z0Z_1_cascade_));
    InMux I__692 (
            .O(N__4078),
            .I(N__4071));
    InMux I__691 (
            .O(N__4077),
            .I(N__4071));
    InMux I__690 (
            .O(N__4076),
            .I(N__4068));
    LocalMux I__689 (
            .O(N__4071),
            .I(countZ0Z_2));
    LocalMux I__688 (
            .O(N__4068),
            .I(countZ0Z_2));
    CascadeMux I__687 (
            .O(N__4063),
            .I(CLKOS3_3_cascade_));
    CascadeMux I__686 (
            .O(N__4060),
            .I(N__4057));
    InMux I__685 (
            .O(N__4057),
            .I(N__4047));
    InMux I__684 (
            .O(N__4056),
            .I(N__4047));
    InMux I__683 (
            .O(N__4055),
            .I(N__4047));
    InMux I__682 (
            .O(N__4054),
            .I(N__4044));
    LocalMux I__681 (
            .O(N__4047),
            .I(countZ0Z_1));
    LocalMux I__680 (
            .O(N__4044),
            .I(countZ0Z_1));
    InMux I__679 (
            .O(N__4039),
            .I(N__4028));
    InMux I__678 (
            .O(N__4038),
            .I(N__4028));
    InMux I__677 (
            .O(N__4037),
            .I(N__4028));
    InMux I__676 (
            .O(N__4036),
            .I(N__4025));
    InMux I__675 (
            .O(N__4035),
            .I(N__4022));
    LocalMux I__674 (
            .O(N__4028),
            .I(countZ0Z_0));
    LocalMux I__673 (
            .O(N__4025),
            .I(countZ0Z_0));
    LocalMux I__672 (
            .O(N__4022),
            .I(countZ0Z_0));
    InMux I__671 (
            .O(N__4015),
            .I(N__4012));
    LocalMux I__670 (
            .O(N__4012),
            .I(G_7_a0_1));
    CascadeMux I__669 (
            .O(N__4009),
            .I(N__4005));
    InMux I__668 (
            .O(N__4008),
            .I(N__4002));
    InMux I__667 (
            .O(N__4005),
            .I(N__3999));
    LocalMux I__666 (
            .O(N__4002),
            .I(count_i_3));
    LocalMux I__665 (
            .O(N__3999),
            .I(count_i_3));
    CascadeMux I__664 (
            .O(N__3994),
            .I(N__3991));
    InMux I__663 (
            .O(N__3991),
            .I(N__3983));
    InMux I__662 (
            .O(N__3990),
            .I(N__3983));
    InMux I__661 (
            .O(N__3989),
            .I(N__3978));
    InMux I__660 (
            .O(N__3988),
            .I(N__3978));
    LocalMux I__659 (
            .O(N__3983),
            .I(CLKOS_i));
    LocalMux I__658 (
            .O(N__3978),
            .I(CLKOS_i));
    InMux I__657 (
            .O(N__3973),
            .I(N__3970));
    LocalMux I__656 (
            .O(N__3970),
            .I(G_7_a0_0));
    CascadeMux I__655 (
            .O(N__3967),
            .I(N__3964));
    InMux I__654 (
            .O(N__3964),
            .I(N__3959));
    InMux I__653 (
            .O(N__3963),
            .I(N__3954));
    InMux I__652 (
            .O(N__3962),
            .I(N__3954));
    LocalMux I__651 (
            .O(N__3959),
            .I(clk_countZ0Z_1));
    LocalMux I__650 (
            .O(N__3954),
            .I(clk_countZ0Z_1));
    CascadeMux I__649 (
            .O(N__3949),
            .I(\uut1.N_217_0_4_cascade_ ));
    CascadeMux I__648 (
            .O(N__3946),
            .I(\uut1.N_216_0_cascade_ ));
    InMux I__647 (
            .O(N__3943),
            .I(N__3939));
    InMux I__646 (
            .O(N__3942),
            .I(N__3936));
    LocalMux I__645 (
            .O(N__3939),
            .I(count_ext_RNIEM1QZ0Z_1));
    LocalMux I__644 (
            .O(N__3936),
            .I(count_ext_RNIEM1QZ0Z_1));
    InMux I__643 (
            .O(N__3931),
            .I(N__3924));
    InMux I__642 (
            .O(N__3930),
            .I(N__3921));
    InMux I__641 (
            .O(N__3929),
            .I(N__3916));
    InMux I__640 (
            .O(N__3928),
            .I(N__3916));
    InMux I__639 (
            .O(N__3927),
            .I(N__3913));
    LocalMux I__638 (
            .O(N__3924),
            .I(count_ext13));
    LocalMux I__637 (
            .O(N__3921),
            .I(count_ext13));
    LocalMux I__636 (
            .O(N__3916),
            .I(count_ext13));
    LocalMux I__635 (
            .O(N__3913),
            .I(count_ext13));
    CascadeMux I__634 (
            .O(N__3904),
            .I(N__3901));
    InMux I__633 (
            .O(N__3901),
            .I(N__3898));
    LocalMux I__632 (
            .O(N__3898),
            .I(N__3894));
    CascadeMux I__631 (
            .O(N__3897),
            .I(N__3890));
    Span4Mux_h I__630 (
            .O(N__3894),
            .I(N__3887));
    InMux I__629 (
            .O(N__3893),
            .I(N__3884));
    InMux I__628 (
            .O(N__3890),
            .I(N__3881));
    Odrv4 I__627 (
            .O(N__3887),
            .I(count_extZ0Z_0));
    LocalMux I__626 (
            .O(N__3884),
            .I(count_extZ0Z_0));
    LocalMux I__625 (
            .O(N__3881),
            .I(count_extZ0Z_0));
    CEMux I__624 (
            .O(N__3874),
            .I(N__3850));
    CEMux I__623 (
            .O(N__3873),
            .I(N__3850));
    CEMux I__622 (
            .O(N__3872),
            .I(N__3850));
    CEMux I__621 (
            .O(N__3871),
            .I(N__3850));
    CEMux I__620 (
            .O(N__3870),
            .I(N__3850));
    CEMux I__619 (
            .O(N__3869),
            .I(N__3850));
    CEMux I__618 (
            .O(N__3868),
            .I(N__3850));
    CEMux I__617 (
            .O(N__3867),
            .I(N__3850));
    GlobalMux I__616 (
            .O(N__3850),
            .I(N__3847));
    gio2CtrlBuf I__615 (
            .O(N__3847),
            .I(N_95_g));
    IoInMux I__614 (
            .O(N__3844),
            .I(N__3841));
    LocalMux I__613 (
            .O(N__3841),
            .I(N__3834));
    InMux I__612 (
            .O(N__3840),
            .I(N__3825));
    InMux I__611 (
            .O(N__3839),
            .I(N__3825));
    InMux I__610 (
            .O(N__3838),
            .I(N__3825));
    InMux I__609 (
            .O(N__3837),
            .I(N__3825));
    IoSpan4Mux I__608 (
            .O(N__3834),
            .I(N__3822));
    LocalMux I__607 (
            .O(N__3825),
            .I(CLKOS_RNI7KOJZ0Z1));
    Odrv4 I__606 (
            .O(N__3822),
            .I(CLKOS_RNI7KOJZ0Z1));
    InMux I__605 (
            .O(N__3817),
            .I(N__3813));
    IoInMux I__604 (
            .O(N__3816),
            .I(N__3810));
    LocalMux I__603 (
            .O(N__3813),
            .I(N__3807));
    LocalMux I__602 (
            .O(N__3810),
            .I(N__3804));
    Span4Mux_s2_v I__601 (
            .O(N__3807),
            .I(N__3800));
    IoSpan4Mux I__600 (
            .O(N__3804),
            .I(N__3797));
    InMux I__599 (
            .O(N__3803),
            .I(N__3794));
    Sp12to4 I__598 (
            .O(N__3800),
            .I(N__3791));
    Span4Mux_s0_v I__597 (
            .O(N__3797),
            .I(N__3786));
    LocalMux I__596 (
            .O(N__3794),
            .I(N__3786));
    Span12Mux_s11_h I__595 (
            .O(N__3791),
            .I(N__3783));
    Sp12to4 I__594 (
            .O(N__3786),
            .I(N__3780));
    Span12Mux_v I__593 (
            .O(N__3783),
            .I(N__3777));
    Span12Mux_v I__592 (
            .O(N__3780),
            .I(N__3774));
    Odrv12 I__591 (
            .O(N__3777),
            .I(test2_c));
    Odrv12 I__590 (
            .O(N__3774),
            .I(test2_c));
    CascadeMux I__589 (
            .O(N__3769),
            .I(N__3764));
    InMux I__588 (
            .O(N__3768),
            .I(N__3761));
    InMux I__587 (
            .O(N__3767),
            .I(N__3758));
    InMux I__586 (
            .O(N__3764),
            .I(N__3755));
    LocalMux I__585 (
            .O(N__3761),
            .I(count_extZ0Z_4));
    LocalMux I__584 (
            .O(N__3758),
            .I(count_extZ0Z_4));
    LocalMux I__583 (
            .O(N__3755),
            .I(count_extZ0Z_4));
    CascadeMux I__582 (
            .O(N__3748),
            .I(\uut1.rx_data_35_0_0_6_cascade_ ));
    CascadeMux I__581 (
            .O(N__3745),
            .I(\uut1.N_218_0_cascade_ ));
    InMux I__580 (
            .O(N__3742),
            .I(N__3739));
    LocalMux I__579 (
            .O(N__3739),
            .I(from_ir_regZ0Z2));
    InMux I__578 (
            .O(N__3736),
            .I(N__3732));
    InMux I__577 (
            .O(N__3735),
            .I(N__3729));
    LocalMux I__576 (
            .O(N__3732),
            .I(from_ir_regZ0Z1));
    LocalMux I__575 (
            .O(N__3729),
            .I(from_ir_regZ0Z1));
    InMux I__574 (
            .O(N__3724),
            .I(N__3720));
    InMux I__573 (
            .O(N__3723),
            .I(N__3717));
    LocalMux I__572 (
            .O(N__3720),
            .I(rst_countZ0Z_8));
    LocalMux I__571 (
            .O(N__3717),
            .I(rst_countZ0Z_8));
    InMux I__570 (
            .O(N__3712),
            .I(N__3708));
    InMux I__569 (
            .O(N__3711),
            .I(N__3705));
    LocalMux I__568 (
            .O(N__3708),
            .I(rst_countZ0Z_7));
    LocalMux I__567 (
            .O(N__3705),
            .I(rst_countZ0Z_7));
    InMux I__566 (
            .O(N__3700),
            .I(N__3697));
    LocalMux I__565 (
            .O(N__3697),
            .I(un1_rst_countlt9_0));
    IoInMux I__564 (
            .O(N__3694),
            .I(N__3691));
    LocalMux I__563 (
            .O(N__3691),
            .I(N__3687));
    IoInMux I__562 (
            .O(N__3690),
            .I(N__3684));
    IoSpan4Mux I__561 (
            .O(N__3687),
            .I(N__3679));
    LocalMux I__560 (
            .O(N__3684),
            .I(N__3679));
    Span4Mux_s3_v I__559 (
            .O(N__3679),
            .I(N__3676));
    Span4Mux_h I__558 (
            .O(N__3676),
            .I(N__3673));
    Odrv4 I__557 (
            .O(N__3673),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__556 (
            .O(N__3670),
            .I(N__3667));
    InMux I__555 (
            .O(N__3667),
            .I(N__3662));
    InMux I__554 (
            .O(N__3666),
            .I(N__3657));
    InMux I__553 (
            .O(N__3665),
            .I(N__3657));
    LocalMux I__552 (
            .O(N__3662),
            .I(N__3654));
    LocalMux I__551 (
            .O(N__3657),
            .I(rst_countZ0Z_0));
    Odrv4 I__550 (
            .O(N__3654),
            .I(rst_countZ0Z_0));
    InMux I__549 (
            .O(N__3649),
            .I(N__3645));
    InMux I__548 (
            .O(N__3648),
            .I(N__3642));
    LocalMux I__547 (
            .O(N__3645),
            .I(N__3639));
    LocalMux I__546 (
            .O(N__3642),
            .I(rst_countZ0Z_1));
    Odrv4 I__545 (
            .O(N__3639),
            .I(rst_countZ0Z_1));
    InMux I__544 (
            .O(N__3634),
            .I(N__3631));
    LocalMux I__543 (
            .O(N__3631),
            .I(N__3628));
    Glb2LocalMux I__542 (
            .O(N__3628),
            .I(N__3616));
    ClkMux I__541 (
            .O(N__3627),
            .I(N__3616));
    ClkMux I__540 (
            .O(N__3626),
            .I(N__3616));
    ClkMux I__539 (
            .O(N__3625),
            .I(N__3616));
    GlobalMux I__538 (
            .O(N__3616),
            .I(N__3613));
    gio2CtrlBuf I__537 (
            .O(N__3613),
            .I(clk_in_c_g));
    CEMux I__536 (
            .O(N__3610),
            .I(N__3601));
    CEMux I__535 (
            .O(N__3609),
            .I(N__3601));
    CEMux I__534 (
            .O(N__3608),
            .I(N__3601));
    GlobalMux I__533 (
            .O(N__3601),
            .I(N__3598));
    gio2CtrlBuf I__532 (
            .O(N__3598),
            .I(un1_rst_countlt21_0_i_g));
    IoInMux I__531 (
            .O(N__3595),
            .I(N__3592));
    LocalMux I__530 (
            .O(N__3592),
            .I(N__3589));
    Odrv12 I__529 (
            .O(N__3589),
            .I(o_rx_data_i_5));
    InMux I__528 (
            .O(N__3586),
            .I(un5_count_ext_cry_1));
    InMux I__527 (
            .O(N__3583),
            .I(un5_count_ext_cry_2));
    InMux I__526 (
            .O(N__3580),
            .I(un5_count_ext_cry_3));
    InMux I__525 (
            .O(N__3577),
            .I(N__3573));
    InMux I__524 (
            .O(N__3576),
            .I(N__3570));
    LocalMux I__523 (
            .O(N__3573),
            .I(count_extZ0Z_3));
    LocalMux I__522 (
            .O(N__3570),
            .I(count_extZ0Z_3));
    InMux I__521 (
            .O(N__3565),
            .I(N__3560));
    InMux I__520 (
            .O(N__3564),
            .I(N__3557));
    InMux I__519 (
            .O(N__3563),
            .I(N__3554));
    LocalMux I__518 (
            .O(N__3560),
            .I(count_extZ0Z_1));
    LocalMux I__517 (
            .O(N__3557),
            .I(count_extZ0Z_1));
    LocalMux I__516 (
            .O(N__3554),
            .I(count_extZ0Z_1));
    InMux I__515 (
            .O(N__3547),
            .I(N__3543));
    InMux I__514 (
            .O(N__3546),
            .I(N__3540));
    LocalMux I__513 (
            .O(N__3543),
            .I(count_extZ0Z_2));
    LocalMux I__512 (
            .O(N__3540),
            .I(count_extZ0Z_2));
    InMux I__511 (
            .O(N__3535),
            .I(N__3531));
    InMux I__510 (
            .O(N__3534),
            .I(N__3528));
    LocalMux I__509 (
            .O(N__3531),
            .I(N__3525));
    LocalMux I__508 (
            .O(N__3528),
            .I(rst_countZ0Z_12));
    Odrv4 I__507 (
            .O(N__3525),
            .I(rst_countZ0Z_12));
    InMux I__506 (
            .O(N__3520),
            .I(rst_count_1_cry_11));
    InMux I__505 (
            .O(N__3517),
            .I(N__3513));
    InMux I__504 (
            .O(N__3516),
            .I(N__3510));
    LocalMux I__503 (
            .O(N__3513),
            .I(N__3507));
    LocalMux I__502 (
            .O(N__3510),
            .I(rst_countZ0Z_13));
    Odrv4 I__501 (
            .O(N__3507),
            .I(rst_countZ0Z_13));
    InMux I__500 (
            .O(N__3502),
            .I(rst_count_1_cry_12));
    InMux I__499 (
            .O(N__3499),
            .I(N__3495));
    InMux I__498 (
            .O(N__3498),
            .I(N__3492));
    LocalMux I__497 (
            .O(N__3495),
            .I(N__3489));
    LocalMux I__496 (
            .O(N__3492),
            .I(rst_countZ0Z_14));
    Odrv4 I__495 (
            .O(N__3489),
            .I(rst_countZ0Z_14));
    InMux I__494 (
            .O(N__3484),
            .I(rst_count_1_cry_13));
    InMux I__493 (
            .O(N__3481),
            .I(N__3477));
    InMux I__492 (
            .O(N__3480),
            .I(N__3474));
    LocalMux I__491 (
            .O(N__3477),
            .I(rst_countZ0Z_15));
    LocalMux I__490 (
            .O(N__3474),
            .I(rst_countZ0Z_15));
    InMux I__489 (
            .O(N__3469),
            .I(rst_count_1_cry_14));
    CascadeMux I__488 (
            .O(N__3466),
            .I(N__3462));
    InMux I__487 (
            .O(N__3465),
            .I(N__3459));
    InMux I__486 (
            .O(N__3462),
            .I(N__3456));
    LocalMux I__485 (
            .O(N__3459),
            .I(rst_countZ0Z_16));
    LocalMux I__484 (
            .O(N__3456),
            .I(rst_countZ0Z_16));
    InMux I__483 (
            .O(N__3451),
            .I(rst_count_1_cry_15));
    InMux I__482 (
            .O(N__3448),
            .I(N__3444));
    InMux I__481 (
            .O(N__3447),
            .I(N__3441));
    LocalMux I__480 (
            .O(N__3444),
            .I(N__3438));
    LocalMux I__479 (
            .O(N__3441),
            .I(rst_countZ0Z_17));
    Odrv4 I__478 (
            .O(N__3438),
            .I(rst_countZ0Z_17));
    InMux I__477 (
            .O(N__3433),
            .I(bfn_6_5_0_));
    InMux I__476 (
            .O(N__3430),
            .I(N__3426));
    InMux I__475 (
            .O(N__3429),
            .I(N__3423));
    LocalMux I__474 (
            .O(N__3426),
            .I(rst_countZ0Z_18));
    LocalMux I__473 (
            .O(N__3423),
            .I(rst_countZ0Z_18));
    InMux I__472 (
            .O(N__3418),
            .I(rst_count_1_cry_17));
    InMux I__471 (
            .O(N__3415),
            .I(N__3412));
    LocalMux I__470 (
            .O(N__3412),
            .I(N__3408));
    CascadeMux I__469 (
            .O(N__3411),
            .I(N__3404));
    Span4Mux_v I__468 (
            .O(N__3408),
            .I(N__3401));
    InMux I__467 (
            .O(N__3407),
            .I(N__3398));
    InMux I__466 (
            .O(N__3404),
            .I(N__3395));
    Odrv4 I__465 (
            .O(N__3401),
            .I(rst_countZ0Z_19));
    LocalMux I__464 (
            .O(N__3398),
            .I(rst_countZ0Z_19));
    LocalMux I__463 (
            .O(N__3395),
            .I(rst_countZ0Z_19));
    InMux I__462 (
            .O(N__3388),
            .I(rst_count_1_cry_18));
    InMux I__461 (
            .O(N__3385),
            .I(rst_count_1_cry_19));
    InMux I__460 (
            .O(N__3382),
            .I(N__3378));
    InMux I__459 (
            .O(N__3381),
            .I(N__3375));
    LocalMux I__458 (
            .O(N__3378),
            .I(rst_countZ0Z_20));
    LocalMux I__457 (
            .O(N__3375),
            .I(rst_countZ0Z_20));
    InMux I__456 (
            .O(N__3370),
            .I(N__3367));
    LocalMux I__455 (
            .O(N__3367),
            .I(rst_countZ0Z_4));
    InMux I__454 (
            .O(N__3364),
            .I(rst_count_1_cry_3));
    InMux I__453 (
            .O(N__3361),
            .I(N__3358));
    LocalMux I__452 (
            .O(N__3358),
            .I(rst_countZ0Z_5));
    InMux I__451 (
            .O(N__3355),
            .I(rst_count_1_cry_4));
    InMux I__450 (
            .O(N__3352),
            .I(N__3349));
    LocalMux I__449 (
            .O(N__3349),
            .I(rst_countZ0Z_6));
    InMux I__448 (
            .O(N__3346),
            .I(rst_count_1_cry_5));
    InMux I__447 (
            .O(N__3343),
            .I(rst_count_1_cry_6));
    InMux I__446 (
            .O(N__3340),
            .I(rst_count_1_cry_7));
    InMux I__445 (
            .O(N__3337),
            .I(N__3333));
    InMux I__444 (
            .O(N__3336),
            .I(N__3330));
    LocalMux I__443 (
            .O(N__3333),
            .I(N__3327));
    LocalMux I__442 (
            .O(N__3330),
            .I(rst_countZ0Z_9));
    Odrv4 I__441 (
            .O(N__3327),
            .I(rst_countZ0Z_9));
    InMux I__440 (
            .O(N__3322),
            .I(bfn_6_4_0_));
    InMux I__439 (
            .O(N__3319),
            .I(N__3315));
    InMux I__438 (
            .O(N__3318),
            .I(N__3312));
    LocalMux I__437 (
            .O(N__3315),
            .I(N__3309));
    LocalMux I__436 (
            .O(N__3312),
            .I(rst_countZ0Z_10));
    Odrv4 I__435 (
            .O(N__3309),
            .I(rst_countZ0Z_10));
    InMux I__434 (
            .O(N__3304),
            .I(rst_count_1_cry_9));
    CascadeMux I__433 (
            .O(N__3301),
            .I(N__3298));
    InMux I__432 (
            .O(N__3298),
            .I(N__3294));
    InMux I__431 (
            .O(N__3297),
            .I(N__3291));
    LocalMux I__430 (
            .O(N__3294),
            .I(N__3288));
    LocalMux I__429 (
            .O(N__3291),
            .I(rst_countZ0Z_11));
    Odrv4 I__428 (
            .O(N__3288),
            .I(rst_countZ0Z_11));
    InMux I__427 (
            .O(N__3283),
            .I(rst_count_1_cry_10));
    InMux I__426 (
            .O(N__3280),
            .I(N__3274));
    InMux I__425 (
            .O(N__3279),
            .I(N__3274));
    LocalMux I__424 (
            .O(N__3274),
            .I(shift_reg2Z0Z_2));
    InMux I__423 (
            .O(N__3271),
            .I(N__3267));
    InMux I__422 (
            .O(N__3270),
            .I(N__3264));
    LocalMux I__421 (
            .O(N__3267),
            .I(shift_reg2Z0Z_3));
    LocalMux I__420 (
            .O(N__3264),
            .I(shift_reg2Z0Z_3));
    CascadeMux I__419 (
            .O(N__3259),
            .I(un1_rst_countlt14_0_cascade_));
    InMux I__418 (
            .O(N__3256),
            .I(N__3253));
    LocalMux I__417 (
            .O(N__3253),
            .I(un1_rst_countlt17));
    InMux I__416 (
            .O(N__3250),
            .I(N__3247));
    LocalMux I__415 (
            .O(N__3247),
            .I(rst_countZ0Z_2));
    InMux I__414 (
            .O(N__3244),
            .I(rst_count_1_cry_1));
    InMux I__413 (
            .O(N__3241),
            .I(N__3238));
    LocalMux I__412 (
            .O(N__3238),
            .I(rst_countZ0Z_3));
    InMux I__411 (
            .O(N__3235),
            .I(rst_count_1_cry_2));
    CascadeMux I__410 (
            .O(N__3232),
            .I(N__3228));
    InMux I__409 (
            .O(N__3231),
            .I(N__3225));
    InMux I__408 (
            .O(N__3228),
            .I(N__3222));
    LocalMux I__407 (
            .O(N__3225),
            .I(shift_reg1Z0Z_3));
    LocalMux I__406 (
            .O(N__3222),
            .I(shift_reg1Z0Z_3));
    InMux I__405 (
            .O(N__3217),
            .I(N__3211));
    InMux I__404 (
            .O(N__3216),
            .I(N__3211));
    LocalMux I__403 (
            .O(N__3211),
            .I(shift_reg1Z0Z_4));
    InMux I__402 (
            .O(N__3208),
            .I(N__3205));
    LocalMux I__401 (
            .O(N__3205),
            .I(un1_rst_countlt18_0));
    IoInMux I__400 (
            .O(N__3202),
            .I(N__3199));
    LocalMux I__399 (
            .O(N__3199),
            .I(N__3196));
    IoSpan4Mux I__398 (
            .O(N__3196),
            .I(N__3193));
    Span4Mux_s0_h I__397 (
            .O(N__3193),
            .I(N__3190));
    Span4Mux_h I__396 (
            .O(N__3190),
            .I(N__3187));
    Odrv4 I__395 (
            .O(N__3187),
            .I(un1_rst_countlt21_0_i));
    InMux I__394 (
            .O(N__3184),
            .I(N__3178));
    InMux I__393 (
            .O(N__3183),
            .I(N__3178));
    LocalMux I__392 (
            .O(N__3178),
            .I(shift_reg2Z0Z_17));
    InMux I__391 (
            .O(N__3175),
            .I(N__3169));
    InMux I__390 (
            .O(N__3174),
            .I(N__3169));
    LocalMux I__389 (
            .O(N__3169),
            .I(shift_reg2Z0Z_16));
    InMux I__388 (
            .O(N__3166),
            .I(N__3162));
    CascadeMux I__387 (
            .O(N__3165),
            .I(N__3159));
    LocalMux I__386 (
            .O(N__3162),
            .I(N__3156));
    InMux I__385 (
            .O(N__3159),
            .I(N__3153));
    Odrv4 I__384 (
            .O(N__3156),
            .I(shift_reg2Z0Z_18));
    LocalMux I__383 (
            .O(N__3153),
            .I(shift_reg2Z0Z_18));
    InMux I__382 (
            .O(N__3148),
            .I(N__3142));
    InMux I__381 (
            .O(N__3147),
            .I(N__3142));
    LocalMux I__380 (
            .O(N__3142),
            .I(shift_reg2Z0Z_0));
    InMux I__379 (
            .O(N__3139),
            .I(N__3136));
    LocalMux I__378 (
            .O(N__3136),
            .I(rx_rdy_13));
    InMux I__377 (
            .O(N__3133),
            .I(N__3130));
    LocalMux I__376 (
            .O(N__3130),
            .I(rx_rdy_5));
    InMux I__375 (
            .O(N__3127),
            .I(N__3121));
    InMux I__374 (
            .O(N__3126),
            .I(N__3121));
    LocalMux I__373 (
            .O(N__3121),
            .I(shift_reg2Z0Z_1));
    InMux I__372 (
            .O(N__3118),
            .I(N__3115));
    LocalMux I__371 (
            .O(N__3115),
            .I(shift_reg1Z0Z_15));
    InMux I__370 (
            .O(N__3112),
            .I(N__3106));
    InMux I__369 (
            .O(N__3111),
            .I(N__3106));
    LocalMux I__368 (
            .O(N__3106),
            .I(shift_reg1Z0Z_10));
    CascadeMux I__367 (
            .O(N__3103),
            .I(N__3099));
    InMux I__366 (
            .O(N__3102),
            .I(N__3094));
    InMux I__365 (
            .O(N__3099),
            .I(N__3094));
    LocalMux I__364 (
            .O(N__3094),
            .I(shift_reg1Z0Z_14));
    InMux I__363 (
            .O(N__3091),
            .I(N__3087));
    InMux I__362 (
            .O(N__3090),
            .I(N__3084));
    LocalMux I__361 (
            .O(N__3087),
            .I(shift_reg1Z0Z_13));
    LocalMux I__360 (
            .O(N__3084),
            .I(shift_reg1Z0Z_13));
    InMux I__359 (
            .O(N__3079),
            .I(N__3073));
    InMux I__358 (
            .O(N__3078),
            .I(N__3073));
    LocalMux I__357 (
            .O(N__3073),
            .I(shift_reg1Z0Z_11));
    InMux I__356 (
            .O(N__3070),
            .I(N__3066));
    InMux I__355 (
            .O(N__3069),
            .I(N__3063));
    LocalMux I__354 (
            .O(N__3066),
            .I(shift_reg1Z0Z_12));
    LocalMux I__353 (
            .O(N__3063),
            .I(shift_reg1Z0Z_12));
    CascadeMux I__352 (
            .O(N__3058),
            .I(N__3054));
    InMux I__351 (
            .O(N__3057),
            .I(N__3051));
    InMux I__350 (
            .O(N__3054),
            .I(N__3048));
    LocalMux I__349 (
            .O(N__3051),
            .I(shift_reg1Z0Z_7));
    LocalMux I__348 (
            .O(N__3048),
            .I(shift_reg1Z0Z_7));
    InMux I__347 (
            .O(N__3043),
            .I(N__3040));
    LocalMux I__346 (
            .O(N__3040),
            .I(i_start_tx_11));
    InMux I__345 (
            .O(N__3037),
            .I(N__3034));
    LocalMux I__344 (
            .O(N__3034),
            .I(i_start_tx_9));
    CascadeMux I__343 (
            .O(N__3031),
            .I(i_start_tx_8_cascade_));
    InMux I__342 (
            .O(N__3028),
            .I(N__3025));
    LocalMux I__341 (
            .O(N__3025),
            .I(i_start_tx_10));
    InMux I__340 (
            .O(N__3022),
            .I(N__3016));
    InMux I__339 (
            .O(N__3021),
            .I(N__3016));
    LocalMux I__338 (
            .O(N__3016),
            .I(shift_reg1Z0Z_5));
    InMux I__337 (
            .O(N__3013),
            .I(N__3009));
    InMux I__336 (
            .O(N__3012),
            .I(N__3006));
    LocalMux I__335 (
            .O(N__3009),
            .I(shift_reg1Z0Z_6));
    LocalMux I__334 (
            .O(N__3006),
            .I(shift_reg1Z0Z_6));
    CascadeMux I__333 (
            .O(N__3001),
            .I(N__2997));
    InMux I__332 (
            .O(N__3000),
            .I(N__2994));
    InMux I__331 (
            .O(N__2997),
            .I(N__2991));
    LocalMux I__330 (
            .O(N__2994),
            .I(shift_reg2Z0Z_4));
    LocalMux I__329 (
            .O(N__2991),
            .I(shift_reg2Z0Z_4));
    InMux I__328 (
            .O(N__2986),
            .I(N__2980));
    InMux I__327 (
            .O(N__2985),
            .I(N__2980));
    LocalMux I__326 (
            .O(N__2980),
            .I(shift_reg2Z0Z_5));
    InMux I__325 (
            .O(N__2977),
            .I(N__2971));
    InMux I__324 (
            .O(N__2976),
            .I(N__2971));
    LocalMux I__323 (
            .O(N__2971),
            .I(shift_reg2Z0Z_6));
    InMux I__322 (
            .O(N__2968),
            .I(N__2962));
    InMux I__321 (
            .O(N__2967),
            .I(N__2962));
    LocalMux I__320 (
            .O(N__2962),
            .I(shift_reg2Z0Z_7));
    InMux I__319 (
            .O(N__2959),
            .I(N__2955));
    CascadeMux I__318 (
            .O(N__2958),
            .I(N__2952));
    LocalMux I__317 (
            .O(N__2955),
            .I(N__2949));
    InMux I__316 (
            .O(N__2952),
            .I(N__2946));
    Odrv4 I__315 (
            .O(N__2949),
            .I(shift_reg2Z0Z_8));
    LocalMux I__314 (
            .O(N__2946),
            .I(shift_reg2Z0Z_8));
    IoInMux I__313 (
            .O(N__2941),
            .I(N__2938));
    LocalMux I__312 (
            .O(N__2938),
            .I(N__2935));
    Span4Mux_s3_h I__311 (
            .O(N__2935),
            .I(N__2932));
    Odrv4 I__310 (
            .O(N__2932),
            .I(GB_BUFFER_clk_in_c_g_THRU_CO));
    CascadeMux I__309 (
            .O(N__2929),
            .I(N__2926));
    InMux I__308 (
            .O(N__2926),
            .I(N__2923));
    LocalMux I__307 (
            .O(N__2923),
            .I(shift_reg2Z0Z_19));
    IoInMux I__306 (
            .O(N__2920),
            .I(N__2917));
    LocalMux I__305 (
            .O(N__2917),
            .I(GB_BUFFER_rst_count_i_g_19_THRU_CO));
    CascadeMux I__304 (
            .O(N__2914),
            .I(N__2910));
    InMux I__303 (
            .O(N__2913),
            .I(N__2907));
    InMux I__302 (
            .O(N__2910),
            .I(N__2904));
    LocalMux I__301 (
            .O(N__2907),
            .I(shift_reg1Z0Z_8));
    LocalMux I__300 (
            .O(N__2904),
            .I(shift_reg1Z0Z_8));
    InMux I__299 (
            .O(N__2899),
            .I(N__2893));
    InMux I__298 (
            .O(N__2898),
            .I(N__2893));
    LocalMux I__297 (
            .O(N__2893),
            .I(shift_reg1Z0Z_9));
    InMux I__296 (
            .O(N__2890),
            .I(N__2884));
    InMux I__295 (
            .O(N__2889),
            .I(N__2884));
    LocalMux I__294 (
            .O(N__2884),
            .I(shift_reg2Z0Z_11));
    InMux I__293 (
            .O(N__2881),
            .I(N__2875));
    InMux I__292 (
            .O(N__2880),
            .I(N__2875));
    LocalMux I__291 (
            .O(N__2875),
            .I(shift_reg2Z0Z_10));
    InMux I__290 (
            .O(N__2872),
            .I(N__2868));
    CascadeMux I__289 (
            .O(N__2871),
            .I(N__2865));
    LocalMux I__288 (
            .O(N__2868),
            .I(N__2862));
    InMux I__287 (
            .O(N__2865),
            .I(N__2859));
    Odrv4 I__286 (
            .O(N__2862),
            .I(shift_reg2Z0Z_12));
    LocalMux I__285 (
            .O(N__2859),
            .I(shift_reg2Z0Z_12));
    InMux I__284 (
            .O(N__2854),
            .I(N__2848));
    InMux I__283 (
            .O(N__2853),
            .I(N__2848));
    LocalMux I__282 (
            .O(N__2848),
            .I(shift_reg2Z0Z_9));
    InMux I__281 (
            .O(N__2845),
            .I(N__2839));
    InMux I__280 (
            .O(N__2844),
            .I(N__2839));
    LocalMux I__279 (
            .O(N__2839),
            .I(shift_reg1Z0Z_1));
    InMux I__278 (
            .O(N__2836),
            .I(N__2830));
    InMux I__277 (
            .O(N__2835),
            .I(N__2830));
    LocalMux I__276 (
            .O(N__2830),
            .I(shift_reg1Z0Z_2));
    InMux I__275 (
            .O(N__2827),
            .I(N__2824));
    LocalMux I__274 (
            .O(N__2824),
            .I(N__2821));
    Odrv4 I__273 (
            .O(N__2821),
            .I(rx_rdy_14));
    CascadeMux I__272 (
            .O(N__2818),
            .I(rx_rdy_16_cascade_));
    InMux I__271 (
            .O(N__2815),
            .I(N__2812));
    LocalMux I__270 (
            .O(N__2812),
            .I(rx_rdy_10));
    InMux I__269 (
            .O(N__2809),
            .I(N__2803));
    InMux I__268 (
            .O(N__2808),
            .I(N__2803));
    LocalMux I__267 (
            .O(N__2803),
            .I(shift_reg1Z0Z_0));
    InMux I__266 (
            .O(N__2800),
            .I(N__2797));
    LocalMux I__265 (
            .O(N__2797),
            .I(rx_rdy_11));
    InMux I__264 (
            .O(N__2794),
            .I(N__2791));
    LocalMux I__263 (
            .O(N__2791),
            .I(N__2787));
    InMux I__262 (
            .O(N__2790),
            .I(N__2784));
    Odrv4 I__261 (
            .O(N__2787),
            .I(shift_reg2Z0Z_15));
    LocalMux I__260 (
            .O(N__2784),
            .I(shift_reg2Z0Z_15));
    IoInMux I__259 (
            .O(N__2779),
            .I(N__2776));
    LocalMux I__258 (
            .O(N__2776),
            .I(N__2773));
    IoSpan4Mux I__257 (
            .O(N__2773),
            .I(N__2770));
    Span4Mux_s2_v I__256 (
            .O(N__2770),
            .I(N__2766));
    IoInMux I__255 (
            .O(N__2769),
            .I(N__2763));
    Sp12to4 I__254 (
            .O(N__2766),
            .I(N__2760));
    LocalMux I__253 (
            .O(N__2763),
            .I(N__2757));
    Odrv12 I__252 (
            .O(N__2760),
            .I(test1_c));
    Odrv4 I__251 (
            .O(N__2757),
            .I(test1_c));
    IoInMux I__250 (
            .O(N__2752),
            .I(N__2749));
    LocalMux I__249 (
            .O(N__2749),
            .I(N__2746));
    Span4Mux_s1_h I__248 (
            .O(N__2746),
            .I(N__2743));
    Odrv4 I__247 (
            .O(N__2743),
            .I(rst_count_i_19));
    IoInMux I__246 (
            .O(N__2740),
            .I(N__2737));
    LocalMux I__245 (
            .O(N__2737),
            .I(N__2734));
    Span4Mux_s1_h I__244 (
            .O(N__2734),
            .I(N__2731));
    Odrv4 I__243 (
            .O(N__2731),
            .I(o_rx_data_i_6));
    InMux I__242 (
            .O(N__2728),
            .I(N__2722));
    InMux I__241 (
            .O(N__2727),
            .I(N__2722));
    LocalMux I__240 (
            .O(N__2722),
            .I(shift_reg2Z0Z_14));
    InMux I__239 (
            .O(N__2719),
            .I(N__2713));
    InMux I__238 (
            .O(N__2718),
            .I(N__2713));
    LocalMux I__237 (
            .O(N__2713),
            .I(shift_reg2Z0Z_13));
    IoInMux I__236 (
            .O(N__2710),
            .I(N__2707));
    LocalMux I__235 (
            .O(N__2707),
            .I(N__2704));
    Span12Mux_s9_v I__234 (
            .O(N__2704),
            .I(N__2701));
    Odrv12 I__233 (
            .O(N__2701),
            .I(\ice_pll_inst.CLKOP ));
    defparam IN_MUX_bfv_7_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_1_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(rst_count_1_cry_8),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(rst_count_1_cry_16),
            .carryinitout(bfn_6_5_0_));
    ICE_GB CLKOS_RNI7KOJ1_0 (
            .USERSIGNALTOGLOBALBUFFER(N__3844),
            .GLOBALBUFFEROUTPUT(N_95_g));
    ICE_GB rst_count_RNIVN0T1_0_20 (
            .USERSIGNALTOGLOBALBUFFER(N__3202),
            .GLOBALBUFFEROUTPUT(un1_rst_countlt21_0_i_g));
    ICE_GB \ice_pll_inst.PLLOUTCORE_derived_clock_RNIPF83  (
            .USERSIGNALTOGLOBALBUFFER(N__2710),
            .GLOBALBUFFEROUTPUT(CLKOP_g));
    ICE_GB count_RNIH42R1_0_2 (
            .USERSIGNALTOGLOBALBUFFER(N__5128),
            .GLOBALBUFFEROUTPUT(N_123_g));
    ICE_GB rst_count_RNI3HF2_0_19 (
            .USERSIGNALTOGLOBALBUFFER(N__2752),
            .GLOBALBUFFEROUTPUT(rst_count_i_g_19));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam rst_count_RNI3HF2_19_LC_2_6_1.C_ON=1'b0;
    defparam rst_count_RNI3HF2_19_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam rst_count_RNI3HF2_19_LC_2_6_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 rst_count_RNI3HF2_19_LC_2_6_1 (
            .in0(N__3415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rst_count_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNISCOA_6_LC_2_7_7 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNISCOA_6_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNISCOA_6_LC_2_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uut1.o_rx_data_RNISCOA_6_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5556),
            .lcout(o_rx_data_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_15_LC_4_1_0.C_ON=1'b0;
    defparam shift_reg2_15_LC_4_1_0.SEQ_MODE=4'b1000;
    defparam shift_reg2_15_LC_4_1_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_15_LC_4_1_0 (
            .in0(N__2728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6044),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_14_LC_4_1_2.C_ON=1'b0;
    defparam shift_reg2_14_LC_4_1_2.SEQ_MODE=4'b1000;
    defparam shift_reg2_14_LC_4_1_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_14_LC_4_1_2 (
            .in0(N__2719),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6044),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_2_0_LC_4_1_5.C_ON=1'b0;
    defparam shift_reg1_RNO_2_0_LC_4_1_5.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_2_0_LC_4_1_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNO_2_0_LC_4_1_5 (
            .in0(N__2790),
            .in1(N__2727),
            .in2(N__2929),
            .in3(N__2718),
            .lcout(rx_rdy_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_13_LC_4_1_7.C_ON=1'b0;
    defparam shift_reg2_13_LC_4_1_7.SEQ_MODE=4'b1000;
    defparam shift_reg2_13_LC_4_1_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_13_LC_4_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2872),
            .lcout(shift_reg2Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6044),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_13_LC_4_2_0.C_ON=1'b0;
    defparam shift_reg1_13_LC_4_2_0.SEQ_MODE=4'b1000;
    defparam shift_reg1_13_LC_4_2_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_13_LC_4_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3070),
            .lcout(shift_reg1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6037),
            .ce(N__3871),
            .sr(_gnd_net_));
    defparam shift_reg1_14_LC_4_2_1.C_ON=1'b0;
    defparam shift_reg1_14_LC_4_2_1.SEQ_MODE=4'b1000;
    defparam shift_reg1_14_LC_4_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_14_LC_4_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3091),
            .lcout(shift_reg1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6037),
            .ce(N__3871),
            .sr(_gnd_net_));
    defparam shift_reg1_7_LC_4_2_2.C_ON=1'b0;
    defparam shift_reg1_7_LC_4_2_2.SEQ_MODE=4'b1000;
    defparam shift_reg1_7_LC_4_2_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_7_LC_4_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3013),
            .lcout(shift_reg1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6037),
            .ce(N__3871),
            .sr(_gnd_net_));
    defparam shift_reg1_8_LC_4_2_6.C_ON=1'b0;
    defparam shift_reg1_8_LC_4_2_6.SEQ_MODE=4'b1000;
    defparam shift_reg1_8_LC_4_2_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_8_LC_4_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3057),
            .lcout(shift_reg1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6037),
            .ce(N__3871),
            .sr(_gnd_net_));
    defparam shift_reg1_9_LC_4_2_7.C_ON=1'b0;
    defparam shift_reg1_9_LC_4_2_7.SEQ_MODE=4'b1000;
    defparam shift_reg1_9_LC_4_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_9_LC_4_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2913),
            .lcout(shift_reg1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6037),
            .ce(N__3871),
            .sr(_gnd_net_));
    defparam shift_reg2_10_LC_4_3_0.C_ON=1'b0;
    defparam shift_reg2_10_LC_4_3_0.SEQ_MODE=4'b1000;
    defparam shift_reg2_10_LC_4_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_10_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2854),
            .lcout(shift_reg2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6031),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_16_LC_4_3_1.C_ON=1'b0;
    defparam shift_reg2_16_LC_4_3_1.SEQ_MODE=4'b1000;
    defparam shift_reg2_16_LC_4_3_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 shift_reg2_16_LC_4_3_1 (
            .in0(_gnd_net_),
            .in1(N__2794),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6031),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_12_LC_4_3_2.C_ON=1'b0;
    defparam shift_reg2_12_LC_4_3_2.SEQ_MODE=4'b1000;
    defparam shift_reg2_12_LC_4_3_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_12_LC_4_3_2 (
            .in0(N__2890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6031),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_9_LC_4_3_4.C_ON=1'b0;
    defparam shift_reg2_9_LC_4_3_4.SEQ_MODE=4'b1000;
    defparam shift_reg2_9_LC_4_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_9_LC_4_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2959),
            .lcout(shift_reg2Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6031),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_11_LC_4_3_5.C_ON=1'b0;
    defparam shift_reg2_11_LC_4_3_5.SEQ_MODE=4'b1000;
    defparam shift_reg2_11_LC_4_3_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_11_LC_4_3_5 (
            .in0(N__2881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6031),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_0_0_LC_4_3_6.C_ON=1'b0;
    defparam shift_reg1_RNO_0_0_LC_4_3_6.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_0_0_LC_4_3_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNO_0_0_LC_4_3_6 (
            .in0(N__2889),
            .in1(N__2880),
            .in2(N__2871),
            .in3(N__2853),
            .lcout(rx_rdy_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNIMSC7_0_LC_4_4_0.C_ON=1'b0;
    defparam shift_reg1_RNIMSC7_0_LC_4_4_0.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNIMSC7_0_LC_4_4_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNIMSC7_0_LC_4_4_0 (
            .in0(N__2808),
            .in1(N__2844),
            .in2(N__3232),
            .in3(N__2835),
            .lcout(i_start_tx_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_1_LC_4_4_1.C_ON=1'b0;
    defparam shift_reg1_1_LC_4_4_1.SEQ_MODE=4'b1000;
    defparam shift_reg1_1_LC_4_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_1_LC_4_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2809),
            .lcout(shift_reg1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6025),
            .ce(N__3874),
            .sr(_gnd_net_));
    defparam shift_reg1_2_LC_4_4_2.C_ON=1'b0;
    defparam shift_reg1_2_LC_4_4_2.SEQ_MODE=4'b1000;
    defparam shift_reg1_2_LC_4_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_2_LC_4_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2845),
            .lcout(shift_reg1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6025),
            .ce(N__3874),
            .sr(_gnd_net_));
    defparam shift_reg1_3_LC_4_4_3.C_ON=1'b0;
    defparam shift_reg1_3_LC_4_4_3.SEQ_MODE=4'b1000;
    defparam shift_reg1_3_LC_4_4_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg1_3_LC_4_4_3 (
            .in0(N__2836),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6025),
            .ce(N__3874),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_3_0_LC_4_4_6.C_ON=1'b0;
    defparam shift_reg1_RNO_3_0_LC_4_4_6.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_3_0_LC_4_4_6.LUT_INIT=16'b0000001000000000;
    LogicCell40 shift_reg1_RNO_3_0_LC_4_4_6 (
            .in0(N__3139),
            .in1(N__3270),
            .in2(N__3001),
            .in3(N__3133),
            .lcout(),
            .ltout(rx_rdy_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_0_LC_4_4_7.C_ON=1'b0;
    defparam shift_reg1_0_LC_4_4_7.SEQ_MODE=4'b1000;
    defparam shift_reg1_0_LC_4_4_7.LUT_INIT=16'b0111111111111111;
    LogicCell40 shift_reg1_0_LC_4_4_7 (
            .in0(N__2827),
            .in1(N__2800),
            .in2(N__2818),
            .in3(N__2815),
            .lcout(shift_reg1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6025),
            .ce(N__3874),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_1_0_LC_4_5_0.C_ON=1'b0;
    defparam shift_reg1_RNO_1_0_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_1_0_LC_4_5_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNO_1_0_LC_4_5_0 (
            .in0(N__2967),
            .in1(N__2976),
            .in2(N__2958),
            .in3(N__2985),
            .lcout(rx_rdy_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_7_LC_4_5_2.C_ON=1'b0;
    defparam shift_reg2_7_LC_4_5_2.SEQ_MODE=4'b1000;
    defparam shift_reg2_7_LC_4_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_7_LC_4_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2977),
            .lcout(shift_reg2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6021),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_5_LC_4_5_3.C_ON=1'b0;
    defparam shift_reg2_5_LC_4_5_3.SEQ_MODE=4'b1000;
    defparam shift_reg2_5_LC_4_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_5_LC_4_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3000),
            .lcout(shift_reg2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6021),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_4_LC_4_5_4.C_ON=1'b0;
    defparam shift_reg2_4_LC_4_5_4.SEQ_MODE=4'b1000;
    defparam shift_reg2_4_LC_4_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_4_LC_4_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3271),
            .lcout(shift_reg2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6021),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_6_LC_4_5_5.C_ON=1'b0;
    defparam shift_reg2_6_LC_4_5_5.SEQ_MODE=4'b1000;
    defparam shift_reg2_6_LC_4_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_6_LC_4_5_5 (
            .in0(N__2986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6021),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_8_LC_4_5_6.C_ON=1'b0;
    defparam shift_reg2_8_LC_4_5_6.SEQ_MODE=4'b1000;
    defparam shift_reg2_8_LC_4_5_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_8_LC_4_5_6 (
            .in0(N__2968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6021),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_in_c_g_THRU_LUT4_0_LC_5_1_0.C_ON=1'b0;
    defparam GB_BUFFER_clk_in_c_g_THRU_LUT4_0_LC_5_1_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_in_c_g_THRU_LUT4_0_LC_5_1_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_in_c_g_THRU_LUT4_0_LC_5_1_0 (
            .in0(N__3634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_in_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_19_LC_5_1_1.C_ON=1'b0;
    defparam shift_reg2_19_LC_5_1_1.SEQ_MODE=4'b1000;
    defparam shift_reg2_19_LC_5_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_19_LC_5_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3166),
            .lcout(shift_reg2Z0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6038),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_rst_count_i_g_19_THRU_LUT4_0_LC_5_1_3.C_ON=1'b0;
    defparam GB_BUFFER_rst_count_i_g_19_THRU_LUT4_0_LC_5_1_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_rst_count_i_g_19_THRU_LUT4_0_LC_5_1_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_rst_count_i_g_19_THRU_LUT4_0_LC_5_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5914),
            .lcout(GB_BUFFER_rst_count_i_g_19_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNI82OT_15_LC_5_2_0.C_ON=1'b0;
    defparam shift_reg1_RNI82OT_15_LC_5_2_0.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNI82OT_15_LC_5_2_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNI82OT_15_LC_5_2_0 (
            .in0(N__3118),
            .in1(N__2898),
            .in2(N__2914),
            .in3(N__3111),
            .lcout(i_start_tx_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_10_LC_5_2_2.C_ON=1'b0;
    defparam shift_reg1_10_LC_5_2_2.SEQ_MODE=4'b1000;
    defparam shift_reg1_10_LC_5_2_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_10_LC_5_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2899),
            .lcout(shift_reg1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6032),
            .ce(N__3869),
            .sr(_gnd_net_));
    defparam shift_reg1_15_LC_5_2_4.C_ON=1'b0;
    defparam shift_reg1_15_LC_5_2_4.SEQ_MODE=4'b1000;
    defparam shift_reg1_15_LC_5_2_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg1_15_LC_5_2_4 (
            .in0(N__3102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6032),
            .ce(N__3869),
            .sr(_gnd_net_));
    defparam shift_reg1_11_LC_5_2_5.C_ON=1'b0;
    defparam shift_reg1_11_LC_5_2_5.SEQ_MODE=4'b1000;
    defparam shift_reg1_11_LC_5_2_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg1_11_LC_5_2_5 (
            .in0(N__3112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6032),
            .ce(N__3869),
            .sr(_gnd_net_));
    defparam shift_reg1_RNIUA2K1_11_LC_5_2_6.C_ON=1'b0;
    defparam shift_reg1_RNIUA2K1_11_LC_5_2_6.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNIUA2K1_11_LC_5_2_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNIUA2K1_11_LC_5_2_6 (
            .in0(N__3078),
            .in1(N__3069),
            .in2(N__3103),
            .in3(N__3090),
            .lcout(i_start_tx_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_12_LC_5_2_7.C_ON=1'b0;
    defparam shift_reg1_12_LC_5_2_7.SEQ_MODE=4'b1000;
    defparam shift_reg1_12_LC_5_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_12_LC_5_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3079),
            .lcout(shift_reg1Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6032),
            .ce(N__3869),
            .sr(_gnd_net_));
    defparam rst_count_RNIVCHL1_15_LC_5_3_0.C_ON=1'b0;
    defparam rst_count_RNIVCHL1_15_LC_5_3_0.SEQ_MODE=4'b0000;
    defparam rst_count_RNIVCHL1_15_LC_5_3_0.LUT_INIT=16'b0000000010000000;
    LogicCell40 rst_count_RNIVCHL1_15_LC_5_3_0 (
            .in0(N__3480),
            .in1(N__3448),
            .in2(N__3466),
            .in3(N__3256),
            .lcout(un1_rst_countlt18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNI6DD7_4_LC_5_3_2.C_ON=1'b0;
    defparam shift_reg1_RNI6DD7_4_LC_5_3_2.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNI6DD7_4_LC_5_3_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNI6DD7_4_LC_5_3_2 (
            .in0(N__3021),
            .in1(N__3012),
            .in2(N__3058),
            .in3(N__3216),
            .lcout(),
            .ltout(i_start_tx_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNI2NK03_0_LC_5_3_3.C_ON=1'b0;
    defparam shift_reg1_RNI2NK03_0_LC_5_3_3.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNI2NK03_0_LC_5_3_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 shift_reg1_RNI2NK03_0_LC_5_3_3 (
            .in0(N__3043),
            .in1(N__3037),
            .in2(N__3031),
            .in3(N__3028),
            .lcout(i_start_tx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_5_LC_5_3_5.C_ON=1'b0;
    defparam shift_reg1_5_LC_5_3_5.SEQ_MODE=4'b1000;
    defparam shift_reg1_5_LC_5_3_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg1_5_LC_5_3_5 (
            .in0(N__3217),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6026),
            .ce(N__3872),
            .sr(_gnd_net_));
    defparam shift_reg1_6_LC_5_3_6.C_ON=1'b0;
    defparam shift_reg1_6_LC_5_3_6.SEQ_MODE=4'b1000;
    defparam shift_reg1_6_LC_5_3_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg1_6_LC_5_3_6 (
            .in0(N__3022),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6026),
            .ce(N__3872),
            .sr(_gnd_net_));
    defparam shift_reg1_4_LC_5_3_7.C_ON=1'b0;
    defparam shift_reg1_4_LC_5_3_7.SEQ_MODE=4'b1000;
    defparam shift_reg1_4_LC_5_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg1_4_LC_5_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3231),
            .lcout(shift_reg1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6026),
            .ce(N__3872),
            .sr(_gnd_net_));
    defparam shift_reg2_18_LC_5_4_0.C_ON=1'b0;
    defparam shift_reg2_18_LC_5_4_0.SEQ_MODE=4'b1000;
    defparam shift_reg2_18_LC_5_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_18_LC_5_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3184),
            .lcout(shift_reg2Z0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6022),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_17_LC_5_4_2.C_ON=1'b0;
    defparam shift_reg2_17_LC_5_4_2.SEQ_MODE=4'b1000;
    defparam shift_reg2_17_LC_5_4_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_17_LC_5_4_2 (
            .in0(N__3175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6022),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_0_LC_5_4_4.C_ON=1'b0;
    defparam shift_reg2_0_LC_5_4_4.SEQ_MODE=4'b1000;
    defparam shift_reg2_0_LC_5_4_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 shift_reg2_0_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__4699),
            .in2(_gnd_net_),
            .in3(N__4717),
            .lcout(shift_reg2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6022),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_1_LC_5_4_5.C_ON=1'b0;
    defparam shift_reg2_1_LC_5_4_5.SEQ_MODE=4'b1000;
    defparam shift_reg2_1_LC_5_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_1_LC_5_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3148),
            .lcout(shift_reg2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6022),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_count_RNIVN0T1_20_LC_5_4_6.C_ON=1'b0;
    defparam rst_count_RNIVN0T1_20_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam rst_count_RNIVN0T1_20_LC_5_4_6.LUT_INIT=16'b0011111101111111;
    LogicCell40 rst_count_RNIVN0T1_20_LC_5_4_6 (
            .in0(N__3208),
            .in1(N__3381),
            .in2(N__3411),
            .in3(N__3429),
            .lcout(un1_rst_countlt21_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_5_0_LC_5_4_7.C_ON=1'b0;
    defparam shift_reg1_RNO_5_0_LC_5_4_7.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_5_0_LC_5_4_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 shift_reg1_RNO_5_0_LC_5_4_7 (
            .in0(N__3183),
            .in1(N__3174),
            .in2(N__3165),
            .in3(N__3147),
            .lcout(rx_rdy_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg1_RNO_4_0_LC_5_5_4.C_ON=1'b0;
    defparam shift_reg1_RNO_4_0_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam shift_reg1_RNO_4_0_LC_5_5_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 shift_reg1_RNO_4_0_LC_5_5_4 (
            .in0(_gnd_net_),
            .in1(N__3279),
            .in2(_gnd_net_),
            .in3(N__3126),
            .lcout(rx_rdy_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_2_LC_5_5_5.C_ON=1'b0;
    defparam shift_reg2_2_LC_5_5_5.SEQ_MODE=4'b1000;
    defparam shift_reg2_2_LC_5_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_reg2_2_LC_5_5_5 (
            .in0(N__3127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_reg2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6018),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_reg2_3_LC_5_5_6.C_ON=1'b0;
    defparam shift_reg2_3_LC_5_5_6.SEQ_MODE=4'b1000;
    defparam shift_reg2_3_LC_5_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_reg2_3_LC_5_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3280),
            .lcout(shift_reg2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6018),
            .ce(),
            .sr(_gnd_net_));
    defparam count_ext_1_LC_6_2_0.C_ON=1'b0;
    defparam count_ext_1_LC_6_2_0.SEQ_MODE=4'b1000;
    defparam count_ext_1_LC_6_2_0.LUT_INIT=16'b0000000000010100;
    LogicCell40 count_ext_1_LC_6_2_0 (
            .in0(N__3943),
            .in1(N__3565),
            .in2(N__3904),
            .in3(N__3931),
            .lcout(count_extZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6024),
            .ce(N__3867),
            .sr(_gnd_net_));
    defparam from_ir_reg2_LC_6_2_4.C_ON=1'b0;
    defparam from_ir_reg2_LC_6_2_4.SEQ_MODE=4'b1000;
    defparam from_ir_reg2_LC_6_2_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 from_ir_reg2_LC_6_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3736),
            .lcout(from_ir_regZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6024),
            .ce(N__3867),
            .sr(_gnd_net_));
    defparam from_ir_reg1_LC_6_2_5.C_ON=1'b0;
    defparam from_ir_reg1_LC_6_2_5.SEQ_MODE=4'b1000;
    defparam from_ir_reg1_LC_6_2_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 from_ir_reg1_LC_6_2_5 (
            .in0(N__3817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(from_ir_regZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6024),
            .ce(N__3867),
            .sr(_gnd_net_));
    defparam rst_count_RNI82L61_10_LC_6_2_6.C_ON=1'b0;
    defparam rst_count_RNI82L61_10_LC_6_2_6.SEQ_MODE=4'b0000;
    defparam rst_count_RNI82L61_10_LC_6_2_6.LUT_INIT=16'b1010000010000000;
    LogicCell40 rst_count_RNI82L61_10_LC_6_2_6 (
            .in0(N__3319),
            .in1(N__3337),
            .in2(N__3301),
            .in3(N__3700),
            .lcout(),
            .ltout(un1_rst_countlt14_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_count_RNIV23E1_12_LC_6_2_7.C_ON=1'b0;
    defparam rst_count_RNIV23E1_12_LC_6_2_7.SEQ_MODE=4'b0000;
    defparam rst_count_RNIV23E1_12_LC_6_2_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 rst_count_RNIV23E1_12_LC_6_2_7 (
            .in0(N__3499),
            .in1(N__3517),
            .in2(N__3259),
            .in3(N__3535),
            .lcout(un1_rst_countlt17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_count_1_cry_1_c_LC_6_3_0.C_ON=1'b1;
    defparam rst_count_1_cry_1_c_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam rst_count_1_cry_1_c_LC_6_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 rst_count_1_cry_1_c_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(N__3649),
            .in2(N__3670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(rst_count_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_count_2_LC_6_3_1.C_ON=1'b1;
    defparam rst_count_2_LC_6_3_1.SEQ_MODE=4'b1000;
    defparam rst_count_2_LC_6_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_2_LC_6_3_1 (
            .in0(_gnd_net_),
            .in1(N__3250),
            .in2(_gnd_net_),
            .in3(N__3244),
            .lcout(rst_countZ0Z_2),
            .ltout(),
            .carryin(rst_count_1_cry_1),
            .carryout(rst_count_1_cry_2),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_3_LC_6_3_2.C_ON=1'b1;
    defparam rst_count_3_LC_6_3_2.SEQ_MODE=4'b1000;
    defparam rst_count_3_LC_6_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_3_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(N__3241),
            .in2(_gnd_net_),
            .in3(N__3235),
            .lcout(rst_countZ0Z_3),
            .ltout(),
            .carryin(rst_count_1_cry_2),
            .carryout(rst_count_1_cry_3),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_4_LC_6_3_3.C_ON=1'b1;
    defparam rst_count_4_LC_6_3_3.SEQ_MODE=4'b1000;
    defparam rst_count_4_LC_6_3_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_4_LC_6_3_3 (
            .in0(_gnd_net_),
            .in1(N__3370),
            .in2(_gnd_net_),
            .in3(N__3364),
            .lcout(rst_countZ0Z_4),
            .ltout(),
            .carryin(rst_count_1_cry_3),
            .carryout(rst_count_1_cry_4),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_5_LC_6_3_4.C_ON=1'b1;
    defparam rst_count_5_LC_6_3_4.SEQ_MODE=4'b1000;
    defparam rst_count_5_LC_6_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_5_LC_6_3_4 (
            .in0(_gnd_net_),
            .in1(N__3361),
            .in2(_gnd_net_),
            .in3(N__3355),
            .lcout(rst_countZ0Z_5),
            .ltout(),
            .carryin(rst_count_1_cry_4),
            .carryout(rst_count_1_cry_5),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_6_LC_6_3_5.C_ON=1'b1;
    defparam rst_count_6_LC_6_3_5.SEQ_MODE=4'b1000;
    defparam rst_count_6_LC_6_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_6_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(N__3352),
            .in2(_gnd_net_),
            .in3(N__3346),
            .lcout(rst_countZ0Z_6),
            .ltout(),
            .carryin(rst_count_1_cry_5),
            .carryout(rst_count_1_cry_6),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_7_LC_6_3_6.C_ON=1'b1;
    defparam rst_count_7_LC_6_3_6.SEQ_MODE=4'b1000;
    defparam rst_count_7_LC_6_3_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_7_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(N__3712),
            .in2(_gnd_net_),
            .in3(N__3343),
            .lcout(rst_countZ0Z_7),
            .ltout(),
            .carryin(rst_count_1_cry_6),
            .carryout(rst_count_1_cry_7),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_8_LC_6_3_7.C_ON=1'b1;
    defparam rst_count_8_LC_6_3_7.SEQ_MODE=4'b1000;
    defparam rst_count_8_LC_6_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_8_LC_6_3_7 (
            .in0(_gnd_net_),
            .in1(N__3724),
            .in2(_gnd_net_),
            .in3(N__3340),
            .lcout(rst_countZ0Z_8),
            .ltout(),
            .carryin(rst_count_1_cry_7),
            .carryout(rst_count_1_cry_8),
            .clk(N__3627),
            .ce(N__3610),
            .sr(_gnd_net_));
    defparam rst_count_9_LC_6_4_0.C_ON=1'b1;
    defparam rst_count_9_LC_6_4_0.SEQ_MODE=4'b1000;
    defparam rst_count_9_LC_6_4_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_9_LC_6_4_0 (
            .in0(_gnd_net_),
            .in1(N__3336),
            .in2(_gnd_net_),
            .in3(N__3322),
            .lcout(rst_countZ0Z_9),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(rst_count_1_cry_9),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_10_LC_6_4_1.C_ON=1'b1;
    defparam rst_count_10_LC_6_4_1.SEQ_MODE=4'b1000;
    defparam rst_count_10_LC_6_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_10_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(N__3318),
            .in2(_gnd_net_),
            .in3(N__3304),
            .lcout(rst_countZ0Z_10),
            .ltout(),
            .carryin(rst_count_1_cry_9),
            .carryout(rst_count_1_cry_10),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_11_LC_6_4_2.C_ON=1'b1;
    defparam rst_count_11_LC_6_4_2.SEQ_MODE=4'b1000;
    defparam rst_count_11_LC_6_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_11_LC_6_4_2 (
            .in0(_gnd_net_),
            .in1(N__3297),
            .in2(_gnd_net_),
            .in3(N__3283),
            .lcout(rst_countZ0Z_11),
            .ltout(),
            .carryin(rst_count_1_cry_10),
            .carryout(rst_count_1_cry_11),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_12_LC_6_4_3.C_ON=1'b1;
    defparam rst_count_12_LC_6_4_3.SEQ_MODE=4'b1000;
    defparam rst_count_12_LC_6_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_12_LC_6_4_3 (
            .in0(_gnd_net_),
            .in1(N__3534),
            .in2(_gnd_net_),
            .in3(N__3520),
            .lcout(rst_countZ0Z_12),
            .ltout(),
            .carryin(rst_count_1_cry_11),
            .carryout(rst_count_1_cry_12),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_13_LC_6_4_4.C_ON=1'b1;
    defparam rst_count_13_LC_6_4_4.SEQ_MODE=4'b1000;
    defparam rst_count_13_LC_6_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_13_LC_6_4_4 (
            .in0(_gnd_net_),
            .in1(N__3516),
            .in2(_gnd_net_),
            .in3(N__3502),
            .lcout(rst_countZ0Z_13),
            .ltout(),
            .carryin(rst_count_1_cry_12),
            .carryout(rst_count_1_cry_13),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_14_LC_6_4_5.C_ON=1'b1;
    defparam rst_count_14_LC_6_4_5.SEQ_MODE=4'b1000;
    defparam rst_count_14_LC_6_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_14_LC_6_4_5 (
            .in0(_gnd_net_),
            .in1(N__3498),
            .in2(_gnd_net_),
            .in3(N__3484),
            .lcout(rst_countZ0Z_14),
            .ltout(),
            .carryin(rst_count_1_cry_13),
            .carryout(rst_count_1_cry_14),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_15_LC_6_4_6.C_ON=1'b1;
    defparam rst_count_15_LC_6_4_6.SEQ_MODE=4'b1000;
    defparam rst_count_15_LC_6_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_15_LC_6_4_6 (
            .in0(_gnd_net_),
            .in1(N__3481),
            .in2(_gnd_net_),
            .in3(N__3469),
            .lcout(rst_countZ0Z_15),
            .ltout(),
            .carryin(rst_count_1_cry_14),
            .carryout(rst_count_1_cry_15),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_16_LC_6_4_7.C_ON=1'b1;
    defparam rst_count_16_LC_6_4_7.SEQ_MODE=4'b1000;
    defparam rst_count_16_LC_6_4_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_16_LC_6_4_7 (
            .in0(_gnd_net_),
            .in1(N__3465),
            .in2(_gnd_net_),
            .in3(N__3451),
            .lcout(rst_countZ0Z_16),
            .ltout(),
            .carryin(rst_count_1_cry_15),
            .carryout(rst_count_1_cry_16),
            .clk(N__3626),
            .ce(N__3609),
            .sr(_gnd_net_));
    defparam rst_count_17_LC_6_5_0.C_ON=1'b1;
    defparam rst_count_17_LC_6_5_0.SEQ_MODE=4'b1000;
    defparam rst_count_17_LC_6_5_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_17_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(N__3447),
            .in2(_gnd_net_),
            .in3(N__3433),
            .lcout(rst_countZ0Z_17),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(rst_count_1_cry_17),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam rst_count_18_LC_6_5_1.C_ON=1'b1;
    defparam rst_count_18_LC_6_5_1.SEQ_MODE=4'b1000;
    defparam rst_count_18_LC_6_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_18_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(N__3430),
            .in2(_gnd_net_),
            .in3(N__3418),
            .lcout(rst_countZ0Z_18),
            .ltout(),
            .carryin(rst_count_1_cry_17),
            .carryout(rst_count_1_cry_18),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam rst_count_19_LC_6_5_2.C_ON=1'b1;
    defparam rst_count_19_LC_6_5_2.SEQ_MODE=4'b1000;
    defparam rst_count_19_LC_6_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 rst_count_19_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(N__3407),
            .in2(_gnd_net_),
            .in3(N__3388),
            .lcout(rst_countZ0Z_19),
            .ltout(),
            .carryin(rst_count_1_cry_18),
            .carryout(rst_count_1_cry_19),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam rst_count_20_LC_6_5_3.C_ON=1'b0;
    defparam rst_count_20_LC_6_5_3.SEQ_MODE=4'b1000;
    defparam rst_count_20_LC_6_5_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 rst_count_20_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(N__3382),
            .in2(_gnd_net_),
            .in3(N__3385),
            .lcout(rst_countZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam rst_count_0_LC_6_5_4.C_ON=1'b0;
    defparam rst_count_0_LC_6_5_4.SEQ_MODE=4'b1000;
    defparam rst_count_0_LC_6_5_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 rst_count_0_LC_6_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3665),
            .lcout(rst_countZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam rst_count_1_LC_6_5_6.C_ON=1'b0;
    defparam rst_count_1_LC_6_5_6.SEQ_MODE=4'b1000;
    defparam rst_count_1_LC_6_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rst_count_1_LC_6_5_6 (
            .in0(_gnd_net_),
            .in1(N__3666),
            .in2(_gnd_net_),
            .in3(N__3648),
            .lcout(rst_countZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3625),
            .ce(N__3608),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNIRBOA_5_LC_6_6_5 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIRBOA_5_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIRBOA_5_LC_6_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uut1.o_rx_data_RNIRBOA_5_LC_6_6_5  (
            .in0(N__5665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_rx_data_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_count_ext_cry_1_c_LC_7_1_0.C_ON=1'b1;
    defparam un5_count_ext_cry_1_c_LC_7_1_0.SEQ_MODE=4'b0000;
    defparam un5_count_ext_cry_1_c_LC_7_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_count_ext_cry_1_c_LC_7_1_0 (
            .in0(_gnd_net_),
            .in1(N__3564),
            .in2(N__3897),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_1_0_),
            .carryout(un5_count_ext_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_ext_2_LC_7_1_1.C_ON=1'b1;
    defparam count_ext_2_LC_7_1_1.SEQ_MODE=4'b1000;
    defparam count_ext_2_LC_7_1_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 count_ext_2_LC_7_1_1 (
            .in0(N__3928),
            .in1(N__3547),
            .in2(_gnd_net_),
            .in3(N__3586),
            .lcout(count_extZ0Z_2),
            .ltout(),
            .carryin(un5_count_ext_cry_1),
            .carryout(un5_count_ext_cry_2),
            .clk(N__6039),
            .ce(N__3868),
            .sr(_gnd_net_));
    defparam count_ext_3_LC_7_1_2.C_ON=1'b1;
    defparam count_ext_3_LC_7_1_2.SEQ_MODE=4'b1000;
    defparam count_ext_3_LC_7_1_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 count_ext_3_LC_7_1_2 (
            .in0(N__3927),
            .in1(N__3577),
            .in2(_gnd_net_),
            .in3(N__3583),
            .lcout(count_extZ0Z_3),
            .ltout(),
            .carryin(un5_count_ext_cry_2),
            .carryout(un5_count_ext_cry_3),
            .clk(N__6039),
            .ce(N__3868),
            .sr(_gnd_net_));
    defparam count_ext_4_LC_7_1_3.C_ON=1'b0;
    defparam count_ext_4_LC_7_1_3.SEQ_MODE=4'b1000;
    defparam count_ext_4_LC_7_1_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 count_ext_4_LC_7_1_3 (
            .in0(N__3929),
            .in1(N__3767),
            .in2(_gnd_net_),
            .in3(N__3580),
            .lcout(count_extZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6039),
            .ce(N__3868),
            .sr(_gnd_net_));
    defparam count_ext_RNIEM1Q_1_LC_7_2_1.C_ON=1'b0;
    defparam count_ext_RNIEM1Q_1_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam count_ext_RNIEM1Q_1_LC_7_2_1.LUT_INIT=16'b0000000000010000;
    LogicCell40 count_ext_RNIEM1Q_1_LC_7_2_1 (
            .in0(N__3576),
            .in1(N__3563),
            .in2(N__3769),
            .in3(N__3546),
            .lcout(count_ext_RNIEM1QZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKOS_RNI7KOJ1_LC_7_2_4.C_ON=1'b0;
    defparam CLKOS_RNI7KOJ1_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam CLKOS_RNI7KOJ1_LC_7_2_4.LUT_INIT=16'b0000000100000000;
    LogicCell40 CLKOS_RNI7KOJ1_LC_7_2_4 (
            .in0(N__4248),
            .in1(N__3990),
            .in2(N__4204),
            .in3(N__4161),
            .lcout(CLKOS_RNI7KOJZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam from_ir_reg2_RNIPD7L_LC_7_2_6.C_ON=1'b0;
    defparam from_ir_reg2_RNIPD7L_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam from_ir_reg2_RNIPD7L_LC_7_2_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 from_ir_reg2_RNIPD7L_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(N__3742),
            .in2(_gnd_net_),
            .in3(N__3735),
            .lcout(count_ext13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKOS_LC_7_2_7.C_ON=1'b0;
    defparam CLKOS_LC_7_2_7.SEQ_MODE=4'b1000;
    defparam CLKOS_LC_7_2_7.LUT_INIT=16'b1111000011010010;
    LogicCell40 CLKOS_LC_7_2_7 (
            .in0(N__4162),
            .in1(N__4202),
            .in2(N__3994),
            .in3(N__4249),
            .lcout(CLKOS_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6033),
            .ce(),
            .sr(_gnd_net_));
    defparam count_3_LC_7_3_0.C_ON=1'b0;
    defparam count_3_LC_7_3_0.SEQ_MODE=4'b1000;
    defparam count_3_LC_7_3_0.LUT_INIT=16'b0111111110000000;
    LogicCell40 count_3_LC_7_3_0 (
            .in0(N__4037),
            .in1(N__4078),
            .in2(N__4060),
            .in3(N__4008),
            .lcout(count_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6027),
            .ce(N__3873),
            .sr(_gnd_net_));
    defparam count_0_LC_7_3_1.C_ON=1'b0;
    defparam count_0_LC_7_3_1.SEQ_MODE=4'b1000;
    defparam count_0_LC_7_3_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 count_0_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4038),
            .lcout(countZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6027),
            .ce(N__3873),
            .sr(_gnd_net_));
    defparam count_2_LC_7_3_2.C_ON=1'b0;
    defparam count_2_LC_7_3_2.SEQ_MODE=4'b1000;
    defparam count_2_LC_7_3_2.LUT_INIT=16'b0111011110001000;
    LogicCell40 count_2_LC_7_3_2 (
            .in0(N__4056),
            .in1(N__4036),
            .in2(_gnd_net_),
            .in3(N__4077),
            .lcout(countZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6027),
            .ce(N__3873),
            .sr(_gnd_net_));
    defparam count_1_LC_7_3_3.C_ON=1'b0;
    defparam count_1_LC_7_3_3.SEQ_MODE=4'b1000;
    defparam count_1_LC_7_3_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 count_1_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(N__4055),
            .in2(_gnd_net_),
            .in3(N__4039),
            .lcout(countZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6027),
            .ce(N__3873),
            .sr(_gnd_net_));
    defparam rst_count_RNI10FM_7_LC_7_3_4.C_ON=1'b0;
    defparam rst_count_RNI10FM_7_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam rst_count_RNI10FM_7_LC_7_3_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 rst_count_RNI10FM_7_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__3723),
            .in2(_gnd_net_),
            .in3(N__3711),
            .lcout(un1_rst_countlt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_4_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_4_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_2_6_LC_7_5_2 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_2_6_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_2_6_LC_7_5_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uut1.rx_data_RNO_2_6_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__4346),
            .in2(_gnd_net_),
            .in3(N__4302),
            .lcout(),
            .ltout(\uut1.rx_data_35_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_6_LC_7_5_3 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_6_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_6_LC_7_5_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uut1.rx_data_RNO_0_6_LC_7_5_3  (
            .in0(N__5191),
            .in1(N__4372),
            .in2(N__3748),
            .in3(N__4931),
            .lcout(),
            .ltout(\uut1.N_218_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_6_LC_7_5_4 .C_ON=1'b0;
    defparam \uut1.rx_data_6_LC_7_5_4 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_6_LC_7_5_4 .LUT_INIT=16'b1110111001001100;
    LogicCell40 \uut1.rx_data_6_LC_7_5_4  (
            .in0(N__4844),
            .in1(N__4642),
            .in2(N__3745),
            .in3(N__4126),
            .lcout(\uut1.rx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6019),
            .ce(),
            .sr(N__5894));
    defparam \uut1.rx_data_7_LC_7_5_6 .C_ON=1'b0;
    defparam \uut1.rx_data_7_LC_7_5_6 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_7_LC_7_5_6 .LUT_INIT=16'b1101100011111000;
    LogicCell40 \uut1.rx_data_7_LC_7_5_6  (
            .in0(N__4845),
            .in1(N__4120),
            .in2(N__4687),
            .in3(N__4090),
            .lcout(\uut1.rx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6019),
            .ce(),
            .sr(N__5894));
    defparam \uut1.state_er_7_LC_7_6_1 .C_ON=1'b0;
    defparam \uut1.state_er_7_LC_7_6_1 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_7_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_7_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4306),
            .lcout(\uut1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_8_LC_7_6_2 .C_ON=1'b0;
    defparam \uut1.state_er_8_LC_7_6_2 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_8_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_8_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4545),
            .lcout(\uut1.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_6_LC_7_6_4 .C_ON=1'b0;
    defparam \uut1.state_er_6_LC_7_6_4 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_6_LC_7_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_6_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4114),
            .lcout(\uut1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_5_LC_7_6_5 .C_ON=1'b0;
    defparam \uut1.state_er_5_LC_7_6_5 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_5_LC_7_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_5_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4352),
            .lcout(\uut1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_4_LC_7_6_6 .C_ON=1'b0;
    defparam \uut1.state_er_4_LC_7_6_6 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_4_LC_7_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_4_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4935),
            .lcout(\uut1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_3_LC_7_6_7 .C_ON=1'b0;
    defparam \uut1.state_er_3_LC_7_6_7 .SEQ_MODE=4'b1010;
    defparam \uut1.state_er_3_LC_7_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.state_er_3_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5189),
            .lcout(\uut1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6016),
            .ce(N__5272),
            .sr(N__5892));
    defparam \uut1.state_er_RNI8D3K1_5_LC_7_7_3 .C_ON=1'b0;
    defparam \uut1.state_er_RNI8D3K1_5_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \uut1.state_er_RNI8D3K1_5_LC_7_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uut1.state_er_RNI8D3K1_5_LC_7_7_3  (
            .in0(N__4928),
            .in1(N__4113),
            .in2(N__4353),
            .in3(N__5179),
            .lcout(\uut1.N_217_0_4 ),
            .ltout(\uut1.N_217_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_3_LC_7_7_4 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_3_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_3_LC_7_7_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uut1.rx_data_RNO_0_3_LC_7_7_4  (
            .in0(N__5007),
            .in1(N__4541),
            .in2(N__3949),
            .in3(N__4303),
            .lcout(\uut1.N_215_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_4_LC_7_7_5 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_4_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_4_LC_7_7_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uut1.rx_data_RNO_0_4_LC_7_7_5  (
            .in0(N__4304),
            .in1(N__4574),
            .in2(N__5018),
            .in3(N__4516),
            .lcout(),
            .ltout(\uut1.N_216_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_4_LC_7_7_6 .C_ON=1'b0;
    defparam \uut1.rx_data_4_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_4_LC_7_7_6 .LUT_INIT=16'b1110111001001100;
    LogicCell40 \uut1.rx_data_4_LC_7_7_6  (
            .in0(N__4843),
            .in1(N__5366),
            .in2(N__3946),
            .in3(N__4381),
            .lcout(\uut1.rx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6015),
            .ce(),
            .sr(N__5891));
    defparam count_ext_0_LC_8_1_0.C_ON=1'b0;
    defparam count_ext_0_LC_8_1_0.SEQ_MODE=4'b1000;
    defparam count_ext_0_LC_8_1_0.LUT_INIT=16'b0000000000010001;
    LogicCell40 count_ext_0_LC_8_1_0 (
            .in0(N__3893),
            .in1(N__3942),
            .in2(_gnd_net_),
            .in3(N__3930),
            .lcout(count_extZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6045),
            .ce(N__3870),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_counter_1_LC_8_2_0 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_1_LC_8_2_0 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_counter_1_LC_8_2_0 .LUT_INIT=16'b0111100001010000;
    LogicCell40 \uut1.rx_sampling_counter_1_LC_8_2_0  (
            .in0(N__3838),
            .in1(N__4402),
            .in2(N__4447),
            .in3(N__4773),
            .lcout(\uut1.rx_sampling_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6040),
            .ce(),
            .sr(N__5904));
    defparam \uut1.rx_sampling_counter_0_LC_8_2_1 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_0_LC_8_2_1 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_counter_0_LC_8_2_1 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \uut1.rx_sampling_counter_0_LC_8_2_1  (
            .in0(N__4401),
            .in1(N__4771),
            .in2(_gnd_net_),
            .in3(N__3837),
            .lcout(\uut1.rx_sampling_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6040),
            .ce(),
            .sr(N__5904));
    defparam \uut1.rx_sampling_counter_3_LC_8_2_2 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_3_LC_8_2_2 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_counter_3_LC_8_2_2 .LUT_INIT=16'b0110110001000100;
    LogicCell40 \uut1.rx_sampling_counter_3_LC_8_2_2  (
            .in0(N__3840),
            .in1(N__4421),
            .in2(N__4483),
            .in3(N__4774),
            .lcout(\uut1.rx_sampling_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6040),
            .ce(),
            .sr(N__5904));
    defparam \uut1.rx_sampling_counter_2_LC_8_2_3 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_2_LC_8_2_3 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_counter_2_LC_8_2_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \uut1.rx_sampling_counter_2_LC_8_2_3  (
            .in0(N__4465),
            .in1(N__4772),
            .in2(N__4474),
            .in3(N__3839),
            .lcout(\uut1.rx_sampling_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6040),
            .ce(),
            .sr(N__5904));
    defparam \uut1.modem_serial_data_LC_8_2_5 .C_ON=1'b0;
    defparam \uut1.modem_serial_data_LC_8_2_5 .SEQ_MODE=4'b1011;
    defparam \uut1.modem_serial_data_LC_8_2_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut1.modem_serial_data_LC_8_2_5  (
            .in0(N__3803),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3768),
            .lcout(\uut1.modem_serial_dataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6040),
            .ce(),
            .sr(N__5904));
    defparam \uut1.rx_sampling_clock_RNO_0_LC_8_3_0 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_RNO_0_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_clock_RNO_0_LC_8_3_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \uut1.rx_sampling_clock_RNO_0_LC_8_3_0  (
            .in0(N__3989),
            .in1(_gnd_net_),
            .in2(N__4247),
            .in3(N__4188),
            .lcout(),
            .ltout(\uut1.rx_sampling_clock_cnv_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_clock_RNO_LC_8_3_1 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_RNO_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_clock_RNO_LC_8_3_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut1.rx_sampling_clock_RNO_LC_8_3_1  (
            .in0(N__4734),
            .in1(N__4972),
            .in2(N__4084),
            .in3(N__4163),
            .lcout(\uut1.rx_sampling_clock_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_RNO_0_1_LC_8_3_2.C_ON=1'b0;
    defparam clk_count_RNO_0_1_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam clk_count_RNO_0_1_LC_8_3_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 clk_count_RNO_0_1_LC_8_3_2 (
            .in0(N__3963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4754),
            .lcout(),
            .ltout(clk_count_RNO_0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_1_LC_8_3_3.C_ON=1'b0;
    defparam clk_count_1_LC_8_3_3.SEQ_MODE=4'b1000;
    defparam clk_count_1_LC_8_3_3.LUT_INIT=16'b1110000011110000;
    LogicCell40 clk_count_1_LC_8_3_3 (
            .in0(N__4189),
            .in1(N__4238),
            .in2(N__4081),
            .in3(N__4164),
            .lcout(clk_countZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6034),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_RNIHMLO_5_LC_8_3_4.C_ON=1'b0;
    defparam clk_count_RNIHMLO_5_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam clk_count_RNIHMLO_5_LC_8_3_4.LUT_INIT=16'b0000000001000000;
    LogicCell40 clk_count_RNIHMLO_5_LC_8_3_4 (
            .in0(N__3962),
            .in1(N__4753),
            .in2(N__4141),
            .in3(N__4260),
            .lcout(CLKOS3_3),
            .ltout(CLKOS3_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIH42R1_2_LC_8_3_5.C_ON=1'b0;
    defparam count_RNIH42R1_2_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam count_RNIH42R1_2_LC_8_3_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 count_RNIH42R1_2_LC_8_3_5 (
            .in0(N__4015),
            .in1(N__4076),
            .in2(N__4063),
            .in3(N__3973),
            .lcout(count_RNIH42R1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNITIVF_1_LC_8_3_6.C_ON=1'b0;
    defparam count_RNITIVF_1_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam count_RNITIVF_1_LC_8_3_6.LUT_INIT=16'b0000000000001000;
    LogicCell40 count_RNITIVF_1_LC_8_3_6 (
            .in0(N__4054),
            .in1(N__4035),
            .in2(N__4246),
            .in3(N__4187),
            .lcout(G_7_a0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIGEIG_3_LC_8_3_7.C_ON=1'b0;
    defparam count_RNIGEIG_3_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam count_RNIGEIG_3_LC_8_3_7.LUT_INIT=16'b0000000000001111;
    LogicCell40 count_RNIGEIG_3_LC_8_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4009),
            .in3(N__3988),
            .lcout(G_7_a0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un3_clk_count_cry_1_c_LC_8_4_0.C_ON=1'b1;
    defparam un3_clk_count_cry_1_c_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un3_clk_count_cry_1_c_LC_8_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un3_clk_count_cry_1_c_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__4755),
            .in2(N__3967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un3_clk_count_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_2_LC_8_4_1.C_ON=1'b1;
    defparam clk_count_2_LC_8_4_1.SEQ_MODE=4'b1000;
    defparam clk_count_2_LC_8_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_count_2_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__4244),
            .in2(_gnd_net_),
            .in3(N__4273),
            .lcout(clk_countZ0Z_2),
            .ltout(),
            .carryin(un3_clk_count_cry_1),
            .carryout(un3_clk_count_cry_2),
            .clk(N__6028),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_RNO_0_3_LC_8_4_2.C_ON=1'b1;
    defparam clk_count_RNO_0_3_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam clk_count_RNO_0_3_LC_8_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_count_RNO_0_3_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__4140),
            .in2(_gnd_net_),
            .in3(N__4270),
            .lcout(clk_count_RNO_0Z0Z_3),
            .ltout(),
            .carryin(un3_clk_count_cry_2),
            .carryout(un3_clk_count_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_4_LC_8_4_3.C_ON=1'b1;
    defparam clk_count_4_LC_8_4_3.SEQ_MODE=4'b1000;
    defparam clk_count_4_LC_8_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_count_4_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(N__4195),
            .in2(_gnd_net_),
            .in3(N__4267),
            .lcout(clk_countZ0Z_4),
            .ltout(),
            .carryin(un3_clk_count_cry_3),
            .carryout(un3_clk_count_cry_4),
            .clk(N__6028),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_5_LC_8_4_4.C_ON=1'b0;
    defparam clk_count_5_LC_8_4_4.SEQ_MODE=4'b1000;
    defparam clk_count_5_LC_8_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_count_5_LC_8_4_4 (
            .in0(_gnd_net_),
            .in1(N__4261),
            .in2(_gnd_net_),
            .in3(N__4264),
            .lcout(clk_countZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6028),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_3_LC_8_4_6.C_ON=1'b0;
    defparam clk_count_3_LC_8_4_6.SEQ_MODE=4'b1000;
    defparam clk_count_3_LC_8_4_6.LUT_INIT=16'b1100100011001100;
    LogicCell40 clk_count_3_LC_8_4_6 (
            .in0(N__4245),
            .in1(N__4210),
            .in2(N__4203),
            .in3(N__4165),
            .lcout(clk_countZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6028),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_6_LC_8_5_0 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_6_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_6_LC_8_5_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \uut1.rx_data_RNO_1_6_LC_8_5_0  (
            .in0(N__4112),
            .in1(N__5318),
            .in2(N__4640),
            .in3(N__5267),
            .lcout(\uut1.rx_data_16_m_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_7_LC_8_5_2 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_7_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_7_LC_8_5_2 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uut1.rx_data_RNO_1_7_LC_8_5_2  (
            .in0(N__5339),
            .in1(N__5268),
            .in2(N__4685),
            .in3(N__4351),
            .lcout(\uut1.rx_data_13_m_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.state_er_RNI3VKT_5_LC_8_5_5 .C_ON=1'b0;
    defparam \uut1.state_er_RNI3VKT_5_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uut1.state_er_RNI3VKT_5_LC_8_5_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uut1.state_er_RNI3VKT_5_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__4301),
            .in2(_gnd_net_),
            .in3(N__4111),
            .lcout(\uut1.N_221_0_2 ),
            .ltout(\uut1.N_221_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_7_LC_8_5_6 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_7_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_7_LC_8_5_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uut1.rx_data_RNO_0_7_LC_8_5_6  (
            .in0(N__4371),
            .in1(N__4930),
            .in2(N__4093),
            .in3(N__5190),
            .lcout(\uut1.N_219_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.state_RNIELAE_1_LC_8_5_7 .C_ON=1'b0;
    defparam \uut1.state_RNIELAE_1_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \uut1.state_RNIELAE_1_LC_8_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uut1.state_RNIELAE_1_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__5340),
            .in2(_gnd_net_),
            .in3(N__5047),
            .lcout(\uut1.state_ns_a2_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_4_LC_8_6_0 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_4_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_4_LC_8_6_0 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \uut1.rx_data_RNO_1_4_LC_8_6_0  (
            .in0(N__5325),
            .in1(N__4540),
            .in2(N__5367),
            .in3(N__5251),
            .lcout(\uut1.rx_data_22_m_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.state_er_RNIV1A91_7_LC_8_6_2 .C_ON=1'b0;
    defparam \uut1.state_er_RNIV1A91_7_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \uut1.state_er_RNIV1A91_7_LC_8_6_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uut1.state_er_RNIV1A91_7_LC_8_6_2  (
            .in0(N__5003),
            .in1(N__4539),
            .in2(_gnd_net_),
            .in3(N__4569),
            .lcout(\uut1.N_221_0_5 ),
            .ltout(\uut1.N_221_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_8_LC_8_6_3 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_8_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_8_LC_8_6_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uut1.rx_data_RNO_0_8_LC_8_6_3  (
            .in0(N__4347),
            .in1(N__5180),
            .in2(N__4375),
            .in3(N__4314),
            .lcout(\uut1.N_220_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_3_LC_8_6_4 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_3_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_3_LC_8_6_4 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uut1.rx_data_RNO_1_3_LC_8_6_4  (
            .in0(N__5324),
            .in1(N__5250),
            .in2(N__4600),
            .in3(N__4570),
            .lcout(\uut1.rx_data_25_m_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_0_9_LC_8_6_5 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_9_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_9_LC_8_6_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uut1.rx_data_RNO_0_9_LC_8_6_5  (
            .in0(N__4370),
            .in1(N__4929),
            .in2(N__4354),
            .in3(N__4315),
            .lcout(\uut1.N_221_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.state_RNID38F_1_LC_8_6_6 .C_ON=1'b0;
    defparam \uut1.state_RNID38F_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \uut1.state_RNID38F_1_LC_8_6_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uut1.state_RNID38F_1_LC_8_6_6  (
            .in0(N__4962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5041),
            .lcout(\uut1.state_RNID38FZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_5_LC_8_6_7 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_5_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_5_LC_8_6_7 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \uut1.rx_data_RNO_1_5_LC_8_6_7  (
            .in0(N__5252),
            .in1(N__5326),
            .in2(N__4804),
            .in3(N__4305),
            .lcout(\uut1.rx_data_19_m_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.state_11_LC_8_7_0 .C_ON=1'b0;
    defparam \uut1.state_11_LC_8_7_0 .SEQ_MODE=4'b1010;
    defparam \uut1.state_11_LC_8_7_0 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \uut1.state_11_LC_8_7_0  (
            .in0(N__4575),
            .in1(N__5446),
            .in2(N__4872),
            .in3(N__5016),
            .lcout(\uut1.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6017),
            .ce(),
            .sr(N__5893));
    defparam \uut1.state_2_LC_8_7_2 .C_ON=1'b0;
    defparam \uut1.state_2_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \uut1.state_2_LC_8_7_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uut1.state_2_LC_8_7_2  (
            .in0(N__4868),
            .in1(N__5447),
            .in2(N__4660),
            .in3(N__5188),
            .lcout(\uut1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6017),
            .ce(),
            .sr(N__5893));
    defparam \uut1.rx_data_3_LC_8_7_4 .C_ON=1'b0;
    defparam \uut1.rx_data_3_LC_8_7_4 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_3_LC_8_7_4 .LUT_INIT=16'b1011100011111000;
    LogicCell40 \uut1.rx_data_3_LC_8_7_4  (
            .in0(N__4618),
            .in1(N__4840),
            .in2(N__4599),
            .in3(N__4612),
            .lcout(\uut1.rx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6017),
            .ce(),
            .sr(N__5893));
    defparam \uut1.rx_data_5_LC_8_7_5 .C_ON=1'b0;
    defparam \uut1.rx_data_5_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_5_LC_8_7_5 .LUT_INIT=16'b1101100011111000;
    LogicCell40 \uut1.rx_data_5_LC_8_7_5  (
            .in0(N__4841),
            .in1(N__4606),
            .in2(N__4803),
            .in3(N__4504),
            .lcout(\uut1.rx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6017),
            .ce(),
            .sr(N__5893));
    defparam \uut1.o_rx_data_6_LC_8_7_7 .C_ON=1'b0;
    defparam \uut1.o_rx_data_6_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_6_LC_8_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut1.o_rx_data_6_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__5422),
            .in2(_gnd_net_),
            .in3(N__4592),
            .lcout(o_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6017),
            .ce(),
            .sr(N__5893));
    defparam \uut1.rx_data_RNO_0_5_LC_8_8_5 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_0_5_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_0_5_LC_8_8_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uut1.rx_data_RNO_0_5_LC_8_8_5  (
            .in0(N__4576),
            .in1(N__4546),
            .in2(N__5017),
            .in3(N__4515),
            .lcout(\uut1.N_217_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_clock_LC_9_2_0 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_LC_9_2_0 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_clock_LC_9_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.rx_sampling_clock_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4422),
            .lcout(\uut1.rx_sampling_clockZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6046),
            .ce(N__4498),
            .sr(N__5907));
    defparam \uut1.rx_sampling_counter_RNO_0_3_LC_9_3_2 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_RNO_0_3_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_counter_RNO_0_3_LC_9_3_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uut1.rx_sampling_counter_RNO_0_3_LC_9_3_2  (
            .in0(N__4400),
            .in1(N__4464),
            .in2(_gnd_net_),
            .in3(N__4443),
            .lcout(\uut1.CO2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_counter_RNO_0_2_LC_9_3_4 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_RNO_0_2_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_counter_RNO_0_2_LC_9_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uut1.rx_sampling_counter_RNO_0_2_LC_9_3_4  (
            .in0(N__4399),
            .in1(N__4463),
            .in2(_gnd_net_),
            .in3(N__4442),
            .lcout(\uut1.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_counter_RNI6JC31_3_LC_9_3_5 .C_ON=1'b0;
    defparam \uut1.rx_sampling_counter_RNI6JC31_3_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_counter_RNI6JC31_3_LC_9_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut1.rx_sampling_counter_RNI6JC31_3_LC_9_3_5  (
            .in0(N__4462),
            .in1(N__4441),
            .in2(N__4423),
            .in3(N__4398),
            .lcout(),
            .ltout(\uut1.rx_sampling_counter16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_sampling_start_RNIQNMM1_LC_9_3_6 .C_ON=1'b0;
    defparam \uut1.rx_sampling_start_RNIQNMM1_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_start_RNIQNMM1_LC_9_3_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \uut1.rx_sampling_start_RNIQNMM1_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(N__4733),
            .in2(N__4777),
            .in3(N__4971),
            .lcout(\uut1.rx_sampling_counter_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_count_0_LC_9_3_7.C_ON=1'b0;
    defparam clk_count_0_LC_9_3_7.SEQ_MODE=4'b1000;
    defparam clk_count_0_LC_9_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_count_0_LC_9_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4756),
            .lcout(clk_countZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6041),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_ready_reg1_LC_9_4_0 .C_ON=1'b0;
    defparam \uut1.rx_data_ready_reg1_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_ready_reg1_LC_9_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.rx_data_ready_reg1_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5413),
            .lcout(\uut1.rx_data_ready_regZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6035),
            .ce(),
            .sr(N__5902));
    defparam \uut1.rx_sampling_start_LC_9_4_5 .C_ON=1'b0;
    defparam \uut1.rx_sampling_start_LC_9_4_5 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_start_LC_9_4_5 .LUT_INIT=16'b0000000000101110;
    LogicCell40 \uut1.rx_sampling_start_LC_9_4_5  (
            .in0(N__4735),
            .in1(N__5046),
            .in2(N__5343),
            .in3(N__4970),
            .lcout(\uut1.rx_sampling_startZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6035),
            .ce(),
            .sr(N__5902));
    defparam \uut1.rx_data_ready_reg2_LC_9_4_6 .C_ON=1'b0;
    defparam \uut1.rx_data_ready_reg2_LC_9_4_6 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_ready_reg2_LC_9_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.rx_data_ready_reg2_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4716),
            .lcout(\uut1.rx_data_ready_regZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6035),
            .ce(),
            .sr(N__5902));
    defparam \uut1.o_rx_data_1_LC_9_5_0 .C_ON=1'b0;
    defparam \uut1.o_rx_data_1_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_1_LC_9_5_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uut1.o_rx_data_1_LC_9_5_0  (
            .in0(N__4888),
            .in1(_gnd_net_),
            .in2(N__5415),
            .in3(_gnd_net_),
            .lcout(o_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.o_rx_data_2_LC_9_5_1 .C_ON=1'b0;
    defparam \uut1.o_rx_data_2_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_2_LC_9_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut1.o_rx_data_2_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__5401),
            .in2(_gnd_net_),
            .in3(N__4686),
            .lcout(o_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.data_validation_LC_9_5_2 .C_ON=1'b0;
    defparam \uut1.data_validation_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \uut1.data_validation_LC_9_5_2 .LUT_INIT=16'b1111110001110000;
    LogicCell40 \uut1.data_validation_LC_9_5_2  (
            .in0(N__4653),
            .in1(N__5261),
            .in2(N__5414),
            .in3(N__5019),
            .lcout(\uut1.data_validationZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.o_rx_data_3_LC_9_5_3 .C_ON=1'b0;
    defparam \uut1.o_rx_data_3_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_3_LC_9_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut1.o_rx_data_3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__5402),
            .in2(_gnd_net_),
            .in3(N__4641),
            .lcout(o_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.state_1_LC_9_5_5 .C_ON=1'b0;
    defparam \uut1.state_1_LC_9_5_5 .SEQ_MODE=4'b1010;
    defparam \uut1.state_1_LC_9_5_5 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \uut1.state_1_LC_9_5_5  (
            .in0(N__5262),
            .in1(N__5045),
            .in2(N__5344),
            .in3(N__4969),
            .lcout(\uut1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.state_0_LC_9_5_6 .C_ON=1'b0;
    defparam \uut1.state_0_LC_9_5_6 .SEQ_MODE=4'b1011;
    defparam \uut1.state_0_LC_9_5_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uut1.state_0_LC_9_5_6  (
            .in0(N__4873),
            .in1(N__5452),
            .in2(_gnd_net_),
            .in3(N__5020),
            .lcout(\uut1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6029),
            .ce(),
            .sr(N__5900));
    defparam \uut1.rx_sampling_clock_reg2_RNIL9O2_LC_9_6_4 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_reg2_RNIL9O2_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_sampling_clock_reg2_RNIL9O2_LC_9_6_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uut1.rx_sampling_clock_reg2_RNIL9O2_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__4864),
            .in2(_gnd_net_),
            .in3(N__5445),
            .lcout(\uut1.rx_sample_en ),
            .ltout(\uut1.rx_sample_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_RNO_1_8_LC_9_6_5 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_8_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_8_LC_9_6_5 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \uut1.rx_data_RNO_1_8_LC_9_6_5  (
            .in0(N__4886),
            .in1(N__5342),
            .in2(N__4939),
            .in3(N__4936),
            .lcout(),
            .ltout(\uut1.rx_data_10_m_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.rx_data_8_LC_9_6_6 .C_ON=1'b0;
    defparam \uut1.rx_data_8_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_8_LC_9_6_6 .LUT_INIT=16'b1110010011101100;
    LogicCell40 \uut1.rx_data_8_LC_9_6_6  (
            .in0(N__4842),
            .in1(N__4887),
            .in2(N__4897),
            .in3(N__4894),
            .lcout(\uut1.rx_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6023),
            .ce(),
            .sr(N__5896));
    defparam \uut1.rx_sampling_clock_reg2_LC_9_7_0 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_reg2_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_clock_reg2_LC_9_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.rx_sampling_clock_reg2_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5451),
            .lcout(\uut1.rx_sampling_clock_regZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.o_rx_data_0_LC_9_7_2 .C_ON=1'b0;
    defparam \uut1.o_rx_data_0_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_0_LC_9_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut1.o_rx_data_0_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__5416),
            .in2(_gnd_net_),
            .in3(N__5210),
            .lcout(o_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.rx_data_9_LC_9_7_4 .C_ON=1'b0;
    defparam \uut1.rx_data_9_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_data_9_LC_9_7_4 .LUT_INIT=16'b1101100011111000;
    LogicCell40 \uut1.rx_data_9_LC_9_7_4  (
            .in0(N__4846),
            .in1(N__5146),
            .in2(N__5217),
            .in3(N__4810),
            .lcout(\uut1.rx_dataZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.o_rx_data_4_LC_9_7_5 .C_ON=1'b0;
    defparam \uut1.o_rx_data_4_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_4_LC_9_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut1.o_rx_data_4_LC_9_7_5  (
            .in0(N__5417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4796),
            .lcout(o_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.rx_sampling_clock_reg1_LC_9_7_6 .C_ON=1'b0;
    defparam \uut1.rx_sampling_clock_reg1_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \uut1.rx_sampling_clock_reg1_LC_9_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut1.rx_sampling_clock_reg1_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5461),
            .lcout(\uut1.rx_sampling_clock_regZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.o_rx_data_5_LC_9_7_7 .C_ON=1'b0;
    defparam \uut1.o_rx_data_5_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \uut1.o_rx_data_5_LC_9_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut1.o_rx_data_5_LC_9_7_7  (
            .in0(N__5418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5368),
            .lcout(o_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6020),
            .ce(),
            .sr(N__5895));
    defparam \uut1.rx_data_RNO_1_9_LC_9_8_0 .C_ON=1'b0;
    defparam \uut1.rx_data_RNO_1_9_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \uut1.rx_data_RNO_1_9_LC_9_8_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \uut1.rx_data_RNO_1_9_LC_9_8_0  (
            .in0(N__5341),
            .in1(N__5266),
            .in2(N__5218),
            .in3(N__5187),
            .lcout(\uut1.rx_data_7_m_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.state_11_LC_11_2_1 .C_ON=1'b0;
    defparam \uut2.state_11_LC_11_2_1 .SEQ_MODE=4'b1010;
    defparam \uut2.state_11_LC_11_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_11_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5140),
            .lcout(\uut2.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6048),
            .ce(N__5938),
            .sr(N__5909));
    defparam \uut2.serial_data_RNO_0_LC_11_3_0 .C_ON=1'b0;
    defparam \uut2.serial_data_RNO_0_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \uut2.serial_data_RNO_0_LC_11_3_0 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \uut2.serial_data_RNO_0_LC_11_3_0  (
            .in0(N__5139),
            .in1(N__5081),
            .in2(N__5127),
            .in3(N__5102),
            .lcout(\uut2.serial_data_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.state_0_LC_11_3_2 .C_ON=1'b0;
    defparam \uut2.state_0_LC_11_3_2 .SEQ_MODE=4'b1011;
    defparam \uut2.state_0_LC_11_3_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uut2.state_0_LC_11_3_2  (
            .in0(N__5527),
            .in1(N__5082),
            .in2(_gnd_net_),
            .in3(N__5104),
            .lcout(\uut2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6047),
            .ce(N__5937),
            .sr(N__5908));
    defparam \uut2.state_13_LC_11_3_3 .C_ON=1'b0;
    defparam \uut2.state_13_LC_11_3_3 .SEQ_MODE=4'b1010;
    defparam \uut2.state_13_LC_11_3_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \uut2.state_13_LC_11_3_3  (
            .in0(N__5103),
            .in1(_gnd_net_),
            .in2(N__5086),
            .in3(_gnd_net_),
            .lcout(\uut2.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6047),
            .ce(N__5937),
            .sr(N__5908));
    defparam \uut2.serial_data_LC_11_4_0 .C_ON=1'b0;
    defparam \uut2.serial_data_LC_11_4_0 .SEQ_MODE=4'b1011;
    defparam \uut2.serial_data_LC_11_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut2.serial_data_LC_11_4_0  (
            .in0(N__5563),
            .in1(N__5497),
            .in2(N__5674),
            .in3(N__5467),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6042),
            .ce(N__5059),
            .sr(N__5905));
    defparam \uut2.serial_data_RNO_3_LC_11_5_0 .C_ON=1'b0;
    defparam \uut2.serial_data_RNO_3_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \uut2.serial_data_RNO_3_LC_11_5_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \uut2.serial_data_RNO_3_LC_11_5_0  (
            .in0(N__5641),
            .in1(N__5598),
            .in2(N__5536),
            .in3(N__6072),
            .lcout(\uut2.serial_data_24_iv_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.tx_data_6_LC_11_6_3 .C_ON=1'b0;
    defparam \uut2.tx_data_6_LC_11_6_3 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_6_LC_11_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_6_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5557),
            .lcout(\uut2.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6030),
            .ce(N__5934),
            .sr(N__5901));
    defparam \uut2.state_10_LC_12_3_0 .C_ON=1'b0;
    defparam \uut2.state_10_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \uut2.state_10_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_10_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5614),
            .lcout(\uut2.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.state_1_LC_12_3_1 .C_ON=1'b0;
    defparam \uut2.state_1_LC_12_3_1 .SEQ_MODE=4'b1010;
    defparam \uut2.state_1_LC_12_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_1_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5491),
            .lcout(\uut2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.state_5_LC_12_3_2 .C_ON=1'b0;
    defparam \uut2.state_5_LC_12_3_2 .SEQ_MODE=4'b1010;
    defparam \uut2.state_5_LC_12_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_5_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5686),
            .lcout(\uut2.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.state_4_LC_12_3_3 .C_ON=1'b0;
    defparam \uut2.state_4_LC_12_3_3 .SEQ_MODE=4'b1010;
    defparam \uut2.state_4_LC_12_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_4_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5479),
            .lcout(\uut2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.state_2_LC_12_3_5 .C_ON=1'b0;
    defparam \uut2.state_2_LC_12_3_5 .SEQ_MODE=4'b1010;
    defparam \uut2.state_2_LC_12_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_2_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5509),
            .lcout(\uut2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.state_3_LC_12_3_7 .C_ON=1'b0;
    defparam \uut2.state_3_LC_12_3_7 .SEQ_MODE=4'b1010;
    defparam \uut2.state_3_LC_12_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_3_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5521),
            .lcout(\uut2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6049),
            .ce(N__5936),
            .sr(N__5910));
    defparam \uut2.serial_data_RNO_2_LC_12_4_1 .C_ON=1'b0;
    defparam \uut2.serial_data_RNO_2_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \uut2.serial_data_RNO_2_LC_12_4_1 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \uut2.serial_data_RNO_2_LC_12_4_1  (
            .in0(N__5626),
            .in1(N__5520),
            .in2(N__5635),
            .in3(N__5508),
            .lcout(\uut2.serial_data_24_iv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.serial_data_RNO_1_LC_12_4_2 .C_ON=1'b0;
    defparam \uut2.serial_data_RNO_1_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \uut2.serial_data_RNO_1_LC_12_4_2 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \uut2.serial_data_RNO_1_LC_12_4_2  (
            .in0(N__5490),
            .in1(N__5610),
            .in2(N__5587),
            .in3(N__5478),
            .lcout(\uut2.serial_data_24_iv_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.serial_data_RNO_4_LC_12_4_5 .C_ON=1'b0;
    defparam \uut2.serial_data_RNO_4_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \uut2.serial_data_RNO_4_LC_12_4_5 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \uut2.serial_data_RNO_4_LC_12_4_5  (
            .in0(N__5620),
            .in1(N__5574),
            .in2(N__6061),
            .in3(N__5685),
            .lcout(\uut2.serial_data_24_iv_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut2.tx_data_5_LC_12_5_0 .C_ON=1'b0;
    defparam \uut2.tx_data_5_LC_12_5_0 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_5_LC_12_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_5_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5664),
            .lcout(\uut2.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.tx_data_1_LC_12_5_1 .C_ON=1'b0;
    defparam \uut2.tx_data_1_LC_12_5_1 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_1_LC_12_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_1_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5775),
            .lcout(\uut2.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.tx_data_0_LC_12_5_2 .C_ON=1'b0;
    defparam \uut2.tx_data_0_LC_12_5_2 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_0_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_0_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5715),
            .lcout(\uut2.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.tx_data_3_LC_12_5_3 .C_ON=1'b0;
    defparam \uut2.tx_data_3_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_3_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_3_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5844),
            .lcout(\uut2.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.state_8_LC_12_5_4 .C_ON=1'b0;
    defparam \uut2.state_8_LC_12_5_4 .SEQ_MODE=4'b1010;
    defparam \uut2.state_8_LC_12_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_8_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5599),
            .lcout(\uut2.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.state_7_LC_12_5_5 .C_ON=1'b0;
    defparam \uut2.state_7_LC_12_5_5 .SEQ_MODE=4'b1010;
    defparam \uut2.state_7_LC_12_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_7_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6073),
            .lcout(\uut2.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.tx_data_2_LC_12_5_6 .C_ON=1'b0;
    defparam \uut2.tx_data_2_LC_12_5_6 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_2_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_2_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5739),
            .lcout(\uut2.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.state_6_LC_12_5_7 .C_ON=1'b0;
    defparam \uut2.state_6_LC_12_5_7 .SEQ_MODE=4'b1010;
    defparam \uut2.state_6_LC_12_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.state_6_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5578),
            .lcout(\uut2.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6043),
            .ce(N__5935),
            .sr(N__5906));
    defparam \uut2.tx_data_4_LC_12_6_6 .C_ON=1'b0;
    defparam \uut2.tx_data_4_LC_12_6_6 .SEQ_MODE=4'b1010;
    defparam \uut2.tx_data_4_LC_12_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut2.tx_data_4_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5812),
            .lcout(\uut2.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6036),
            .ce(N__5933),
            .sr(N__5903));
    defparam \uut1.o_rx_data_RNIP9OA_3_LC_12_7_1 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIP9OA_3_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIP9OA_3_LC_12_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uut1.o_rx_data_RNIP9OA_3_LC_12_7_1  (
            .in0(N__5848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_rx_data_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNIQAOA_4_LC_12_7_4 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIQAOA_4_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIQAOA_4_LC_12_7_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \uut1.o_rx_data_RNIQAOA_4_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__5811),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_rx_data_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNIN7OA_1_LC_12_9_6 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIN7OA_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIN7OA_1_LC_12_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uut1.o_rx_data_RNIN7OA_1_LC_12_9_6  (
            .in0(N__5779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_rx_data_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNIO8OA_2_LC_12_11_3 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIO8OA_2_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIO8OA_2_LC_12_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uut1.o_rx_data_RNIO8OA_2_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5746),
            .lcout(o_rx_data_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut1.o_rx_data_RNIM6OA_0_LC_12_11_4 .C_ON=1'b0;
    defparam \uut1.o_rx_data_RNIM6OA_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \uut1.o_rx_data_RNIM6OA_0_LC_12_11_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \uut1.o_rx_data_RNIM6OA_0_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__5716),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_rx_data_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // uart
